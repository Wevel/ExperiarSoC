magic
tech sky130A
magscale 1 2
timestamp 1654557607
<< viali >>
rect 2329 39593 2363 39627
rect 3065 39593 3099 39627
rect 3985 39593 4019 39627
rect 27169 39593 27203 39627
rect 41429 39593 41463 39627
rect 48973 39593 49007 39627
rect 56425 39593 56459 39627
rect 19257 39457 19291 39491
rect 1409 39389 1443 39423
rect 2145 39389 2179 39423
rect 2881 39389 2915 39423
rect 3801 39389 3835 39423
rect 26985 39389 27019 39423
rect 33793 39389 33827 39423
rect 56241 39389 56275 39423
rect 1593 39253 1627 39287
rect 34069 39253 34103 39287
rect 32137 39049 32171 39083
rect 1409 38913 1443 38947
rect 32321 38913 32355 38947
rect 1593 38709 1627 38743
rect 1593 38505 1627 38539
rect 1409 38301 1443 38335
rect 1409 37825 1443 37859
rect 1593 37621 1627 37655
rect 1409 36737 1443 36771
rect 1593 36601 1627 36635
rect 1409 36125 1443 36159
rect 1593 35989 1627 36023
rect 1869 34969 1903 35003
rect 1961 34901 1995 34935
rect 1593 34697 1627 34731
rect 2145 34697 2179 34731
rect 1409 34561 1443 34595
rect 2329 34561 2363 34595
rect 1409 33949 1443 33983
rect 1593 33813 1627 33847
rect 1409 33473 1443 33507
rect 2513 33473 2547 33507
rect 1685 33405 1719 33439
rect 2329 33269 2363 33303
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 1409 32385 1443 32419
rect 1593 32181 1627 32215
rect 2145 31977 2179 32011
rect 1409 31773 1443 31807
rect 2329 31773 2363 31807
rect 1593 31637 1627 31671
rect 1777 31297 1811 31331
rect 2513 31229 2547 31263
rect 1409 30685 1443 30719
rect 2421 30685 2455 30719
rect 3065 30685 3099 30719
rect 4905 30685 4939 30719
rect 1593 30549 1627 30583
rect 2237 30549 2271 30583
rect 2881 30549 2915 30583
rect 4721 30549 4755 30583
rect 4712 30277 4746 30311
rect 1593 30209 1627 30243
rect 2320 30209 2354 30243
rect 4445 30209 4479 30243
rect 2053 30141 2087 30175
rect 1409 30005 1443 30039
rect 3433 30005 3467 30039
rect 5825 30005 5859 30039
rect 2329 29801 2363 29835
rect 4537 29801 4571 29835
rect 6377 29801 6411 29835
rect 2789 29665 2823 29699
rect 2973 29665 3007 29699
rect 4997 29665 5031 29699
rect 5089 29665 5123 29699
rect 6469 29665 6503 29699
rect 1685 29597 1719 29631
rect 4905 29597 4939 29631
rect 6653 29597 6687 29631
rect 2697 29529 2731 29563
rect 6377 29529 6411 29563
rect 1777 29461 1811 29495
rect 6837 29461 6871 29495
rect 5641 29257 5675 29291
rect 7757 29257 7791 29291
rect 12909 29257 12943 29291
rect 15485 29257 15519 29291
rect 6622 29189 6656 29223
rect 1409 29121 1443 29155
rect 2789 29121 2823 29155
rect 5825 29121 5859 29155
rect 11529 29121 11563 29155
rect 11796 29121 11830 29155
rect 14105 29121 14139 29155
rect 14372 29121 14406 29155
rect 6377 29053 6411 29087
rect 1593 28985 1627 29019
rect 2605 28985 2639 29019
rect 2513 28713 2547 28747
rect 6193 28713 6227 28747
rect 12173 28713 12207 28747
rect 14749 28713 14783 28747
rect 3065 28577 3099 28611
rect 6653 28577 6687 28611
rect 6837 28577 6871 28611
rect 6561 28509 6595 28543
rect 12357 28509 12391 28543
rect 12633 28509 12667 28543
rect 14933 28509 14967 28543
rect 15209 28509 15243 28543
rect 17325 28509 17359 28543
rect 1869 28441 1903 28475
rect 2973 28441 3007 28475
rect 12541 28441 12575 28475
rect 15117 28441 15151 28475
rect 17592 28441 17626 28475
rect 1961 28373 1995 28407
rect 2881 28373 2915 28407
rect 18705 28373 18739 28407
rect 17049 28169 17083 28203
rect 18061 28169 18095 28203
rect 2780 28101 2814 28135
rect 18429 28101 18463 28135
rect 1409 28033 1443 28067
rect 16865 28033 16899 28067
rect 17141 28033 17175 28067
rect 18245 28033 18279 28067
rect 18521 28033 18555 28067
rect 2513 27965 2547 27999
rect 3893 27897 3927 27931
rect 1593 27829 1627 27863
rect 16681 27829 16715 27863
rect 16681 27625 16715 27659
rect 2145 27489 2179 27523
rect 15301 27489 15335 27523
rect 2881 27421 2915 27455
rect 3985 27421 4019 27455
rect 5365 27421 5399 27455
rect 5825 27421 5859 27455
rect 10149 27421 10183 27455
rect 15568 27421 15602 27455
rect 1869 27353 1903 27387
rect 6070 27353 6104 27387
rect 10416 27353 10450 27387
rect 2697 27285 2731 27319
rect 3801 27285 3835 27319
rect 5181 27285 5215 27319
rect 7205 27285 7239 27319
rect 11529 27285 11563 27319
rect 6377 27081 6411 27115
rect 6837 27081 6871 27115
rect 9597 27081 9631 27115
rect 10517 27081 10551 27115
rect 10885 27081 10919 27115
rect 14749 27081 14783 27115
rect 2228 27013 2262 27047
rect 3985 26945 4019 26979
rect 6745 26945 6779 26979
rect 8484 26945 8518 26979
rect 10701 26945 10735 26979
rect 10977 26945 11011 26979
rect 13369 26945 13403 26979
rect 13636 26945 13670 26979
rect 17877 26945 17911 26979
rect 18144 26945 18178 26979
rect 1961 26877 1995 26911
rect 6929 26877 6963 26911
rect 8217 26877 8251 26911
rect 3341 26809 3375 26843
rect 3801 26741 3835 26775
rect 19257 26741 19291 26775
rect 2329 26537 2363 26571
rect 9137 26537 9171 26571
rect 12449 26537 12483 26571
rect 14749 26537 14783 26571
rect 17509 26537 17543 26571
rect 18245 26537 18279 26571
rect 4353 26469 4387 26503
rect 2789 26401 2823 26435
rect 2881 26401 2915 26435
rect 4997 26401 5031 26435
rect 16129 26401 16163 26435
rect 1409 26333 1443 26367
rect 4537 26333 4571 26367
rect 5253 26333 5287 26367
rect 9321 26333 9355 26367
rect 9505 26333 9539 26367
rect 9597 26333 9631 26367
rect 14105 26333 14139 26367
rect 14253 26333 14287 26367
rect 14473 26333 14507 26367
rect 14570 26333 14604 26367
rect 18429 26333 18463 26367
rect 18613 26333 18647 26367
rect 18705 26333 18739 26367
rect 2697 26265 2731 26299
rect 12357 26265 12391 26299
rect 14381 26265 14415 26299
rect 15025 26265 15059 26299
rect 16374 26265 16408 26299
rect 1593 26197 1627 26231
rect 6377 26197 6411 26231
rect 3985 25993 4019 26027
rect 4537 25993 4571 26027
rect 4997 25993 5031 26027
rect 16129 25993 16163 26027
rect 4905 25925 4939 25959
rect 15853 25925 15887 25959
rect 1869 25857 1903 25891
rect 2881 25857 2915 25891
rect 3893 25857 3927 25891
rect 12633 25857 12667 25891
rect 12900 25857 12934 25891
rect 15485 25857 15519 25891
rect 15633 25857 15667 25891
rect 15761 25857 15795 25891
rect 15950 25857 15984 25891
rect 5089 25789 5123 25823
rect 2697 25721 2731 25755
rect 2145 25653 2179 25687
rect 14013 25653 14047 25687
rect 14749 25381 14783 25415
rect 1409 25245 1443 25279
rect 2513 25245 2547 25279
rect 5641 25245 5675 25279
rect 8953 25245 8987 25279
rect 10793 25245 10827 25279
rect 14105 25245 14139 25279
rect 14253 25245 14287 25279
rect 14473 25245 14507 25279
rect 14570 25245 14604 25279
rect 6377 25177 6411 25211
rect 9220 25177 9254 25211
rect 11060 25177 11094 25211
rect 14381 25177 14415 25211
rect 1593 25109 1627 25143
rect 2329 25109 2363 25143
rect 5457 25109 5491 25143
rect 6653 25109 6687 25143
rect 10333 25109 10367 25143
rect 12173 25109 12207 25143
rect 15025 25109 15059 25143
rect 5549 24905 5583 24939
rect 10333 24905 10367 24939
rect 10057 24837 10091 24871
rect 1593 24769 1627 24803
rect 2412 24769 2446 24803
rect 5457 24769 5491 24803
rect 6633 24769 6667 24803
rect 9689 24769 9723 24803
rect 9782 24769 9816 24803
rect 9965 24769 9999 24803
rect 10154 24769 10188 24803
rect 19145 24769 19179 24803
rect 2145 24701 2179 24735
rect 5641 24701 5675 24735
rect 6377 24701 6411 24735
rect 18889 24701 18923 24735
rect 3525 24633 3559 24667
rect 1409 24565 1443 24599
rect 5089 24565 5123 24599
rect 7757 24565 7791 24599
rect 20269 24565 20303 24599
rect 2329 24361 2363 24395
rect 10977 24361 11011 24395
rect 18245 24361 18279 24395
rect 2789 24225 2823 24259
rect 2881 24225 2915 24259
rect 5181 24225 5215 24259
rect 15577 24225 15611 24259
rect 19257 24225 19291 24259
rect 1501 24157 1535 24191
rect 2697 24157 2731 24191
rect 10333 24157 10367 24191
rect 10481 24157 10515 24191
rect 10798 24157 10832 24191
rect 12909 24157 12943 24191
rect 13002 24157 13036 24191
rect 13277 24157 13311 24191
rect 13415 24157 13449 24191
rect 18429 24157 18463 24191
rect 18705 24157 18739 24191
rect 4997 24089 5031 24123
rect 10609 24089 10643 24123
rect 10701 24089 10735 24123
rect 13185 24089 13219 24123
rect 15844 24089 15878 24123
rect 18613 24089 18647 24123
rect 19502 24089 19536 24123
rect 1777 24021 1811 24055
rect 13553 24021 13587 24055
rect 16957 24021 16991 24055
rect 20637 24021 20671 24055
rect 1593 23817 1627 23851
rect 15853 23817 15887 23851
rect 19073 23817 19107 23851
rect 6377 23749 6411 23783
rect 12173 23749 12207 23783
rect 13084 23749 13118 23783
rect 15485 23749 15519 23783
rect 15577 23749 15611 23783
rect 1409 23681 1443 23715
rect 2145 23681 2179 23715
rect 2412 23681 2446 23715
rect 6653 23681 6687 23715
rect 9128 23681 9162 23715
rect 11989 23681 12023 23715
rect 15209 23681 15243 23715
rect 15357 23681 15391 23715
rect 15674 23681 15708 23715
rect 19257 23681 19291 23715
rect 19441 23681 19475 23715
rect 19533 23681 19567 23715
rect 6469 23613 6503 23647
rect 8861 23613 8895 23647
rect 12817 23613 12851 23647
rect 10241 23545 10275 23579
rect 3525 23477 3559 23511
rect 6377 23477 6411 23511
rect 6837 23477 6871 23511
rect 14197 23477 14231 23511
rect 2697 23273 2731 23307
rect 5825 23273 5859 23307
rect 6469 23273 6503 23307
rect 10425 23273 10459 23307
rect 14841 23273 14875 23307
rect 6009 23205 6043 23239
rect 13461 23205 13495 23239
rect 1409 23137 1443 23171
rect 5733 23137 5767 23171
rect 6653 23137 6687 23171
rect 16037 23137 16071 23171
rect 1685 23069 1719 23103
rect 2881 23069 2915 23103
rect 3985 23069 4019 23103
rect 5825 23069 5859 23103
rect 6745 23069 6779 23103
rect 9781 23069 9815 23103
rect 9929 23069 9963 23103
rect 10149 23069 10183 23103
rect 10246 23069 10280 23103
rect 11713 23069 11747 23103
rect 13277 23069 13311 23103
rect 14749 23069 14783 23103
rect 21741 23069 21775 23103
rect 25421 23069 25455 23103
rect 28641 23069 28675 23103
rect 31217 23069 31251 23103
rect 5549 23001 5583 23035
rect 6469 23001 6503 23035
rect 10057 23001 10091 23035
rect 12541 23001 12575 23035
rect 12725 23001 12759 23035
rect 16304 23001 16338 23035
rect 22008 23001 22042 23035
rect 25688 23001 25722 23035
rect 31484 23001 31518 23035
rect 3801 22933 3835 22967
rect 6929 22933 6963 22967
rect 11897 22933 11931 22967
rect 17417 22933 17451 22967
rect 23121 22933 23155 22967
rect 26801 22933 26835 22967
rect 28457 22933 28491 22967
rect 32597 22933 32631 22967
rect 2237 22729 2271 22763
rect 2697 22729 2731 22763
rect 16773 22729 16807 22763
rect 25789 22729 25823 22763
rect 26157 22729 26191 22763
rect 27997 22729 28031 22763
rect 32597 22729 32631 22763
rect 17141 22661 17175 22695
rect 27813 22661 27847 22695
rect 28702 22661 28736 22695
rect 32229 22661 32263 22695
rect 32429 22661 32463 22695
rect 1409 22593 1443 22627
rect 2605 22593 2639 22627
rect 3976 22593 4010 22627
rect 7113 22593 7147 22627
rect 7205 22593 7239 22627
rect 7389 22593 7423 22627
rect 7481 22593 7515 22627
rect 11529 22593 11563 22627
rect 16957 22593 16991 22627
rect 17233 22593 17267 22627
rect 18429 22593 18463 22627
rect 18521 22593 18555 22627
rect 19533 22593 19567 22627
rect 19717 22593 19751 22627
rect 22192 22593 22226 22627
rect 25973 22593 26007 22627
rect 26249 22593 26283 22627
rect 27629 22593 27663 22627
rect 31401 22593 31435 22627
rect 31585 22593 31619 22627
rect 33609 22593 33643 22627
rect 33793 22593 33827 22627
rect 34621 22593 34655 22627
rect 34877 22593 34911 22627
rect 2789 22525 2823 22559
rect 3709 22525 3743 22559
rect 18613 22525 18647 22559
rect 18705 22525 18739 22559
rect 19437 22525 19471 22559
rect 19625 22525 19659 22559
rect 21925 22525 21959 22559
rect 28457 22525 28491 22559
rect 1593 22389 1627 22423
rect 5089 22389 5123 22423
rect 6929 22389 6963 22423
rect 11713 22389 11747 22423
rect 18245 22389 18279 22423
rect 19257 22389 19291 22423
rect 23305 22389 23339 22423
rect 29837 22389 29871 22423
rect 31401 22389 31435 22423
rect 32413 22389 32447 22423
rect 33977 22389 34011 22423
rect 36001 22389 36035 22423
rect 11989 22185 12023 22219
rect 20361 22185 20395 22219
rect 23029 22185 23063 22219
rect 28365 22185 28399 22219
rect 31493 22185 31527 22219
rect 34713 22185 34747 22219
rect 19349 22117 19383 22151
rect 4445 22049 4479 22083
rect 10609 22049 10643 22083
rect 14105 22049 14139 22083
rect 18153 22049 18187 22083
rect 18337 22049 18371 22083
rect 18521 22049 18555 22083
rect 19534 22049 19568 22083
rect 19809 22049 19843 22083
rect 20637 22049 20671 22083
rect 20729 22049 20763 22083
rect 32965 22049 32999 22083
rect 1869 21981 1903 22015
rect 2881 21981 2915 22015
rect 4261 21981 4295 22015
rect 7205 21981 7239 22015
rect 7481 21981 7515 22015
rect 7941 21981 7975 22015
rect 12633 21981 12667 22015
rect 12817 21981 12851 22015
rect 12909 21981 12943 22015
rect 18429 21981 18463 22015
rect 18613 21981 18647 22015
rect 19625 21981 19659 22015
rect 19717 21981 19751 22015
rect 20545 21981 20579 22015
rect 20821 21981 20855 22015
rect 22293 21981 22327 22015
rect 22569 21981 22603 22015
rect 23213 21981 23247 22015
rect 23489 21981 23523 22015
rect 28641 21981 28675 22015
rect 28733 21981 28767 22015
rect 28825 21981 28859 22015
rect 29009 21981 29043 22015
rect 30205 21981 30239 22015
rect 30481 21981 30515 22015
rect 31677 21981 31711 22015
rect 31953 21981 31987 22015
rect 33241 21981 33275 22015
rect 33333 21981 33367 22015
rect 33425 21981 33459 22015
rect 33609 21981 33643 22015
rect 34897 21981 34931 22015
rect 37933 21981 37967 22015
rect 2237 21913 2271 21947
rect 4353 21913 4387 21947
rect 10876 21913 10910 21947
rect 12449 21913 12483 21947
rect 14350 21913 14384 21947
rect 23397 21913 23431 21947
rect 38200 21913 38234 21947
rect 2697 21845 2731 21879
rect 3893 21845 3927 21879
rect 7021 21845 7055 21879
rect 7389 21845 7423 21879
rect 8125 21845 8159 21879
rect 15485 21845 15519 21879
rect 22109 21845 22143 21879
rect 22477 21845 22511 21879
rect 31861 21845 31895 21879
rect 39313 21845 39347 21879
rect 3893 21641 3927 21675
rect 13829 21641 13863 21675
rect 16681 21641 16715 21675
rect 19073 21641 19107 21675
rect 29101 21641 29135 21675
rect 31493 21641 31527 21675
rect 33057 21641 33091 21675
rect 33793 21641 33827 21675
rect 35725 21641 35759 21675
rect 14197 21573 14231 21607
rect 32965 21573 32999 21607
rect 35357 21573 35391 21607
rect 36277 21573 36311 21607
rect 1409 21505 1443 21539
rect 2421 21505 2455 21539
rect 3065 21505 3099 21539
rect 4077 21505 4111 21539
rect 6929 21505 6963 21539
rect 7205 21505 7239 21539
rect 7849 21505 7883 21539
rect 8677 21505 8711 21539
rect 8861 21505 8895 21539
rect 14013 21505 14047 21539
rect 14289 21505 14323 21539
rect 14841 21505 14875 21539
rect 17049 21505 17083 21539
rect 17969 21505 18003 21539
rect 19257 21505 19291 21539
rect 19441 21505 19475 21539
rect 24952 21505 24986 21539
rect 29009 21505 29043 21539
rect 29193 21505 29227 21539
rect 31309 21505 31343 21539
rect 31585 21505 31619 21539
rect 32689 21505 32723 21539
rect 32873 21505 32907 21539
rect 33241 21505 33275 21539
rect 33701 21505 33735 21539
rect 35081 21505 35115 21539
rect 35174 21505 35208 21539
rect 35449 21505 35483 21539
rect 35587 21505 35621 21539
rect 38761 21505 38795 21539
rect 7113 21437 7147 21471
rect 7941 21437 7975 21471
rect 16865 21437 16899 21471
rect 16957 21437 16991 21471
rect 17141 21437 17175 21471
rect 17877 21437 17911 21471
rect 18061 21437 18095 21471
rect 18153 21437 18187 21471
rect 19349 21437 19383 21471
rect 19533 21437 19567 21471
rect 24685 21437 24719 21471
rect 38853 21437 38887 21471
rect 8769 21369 8803 21403
rect 15025 21369 15059 21403
rect 31309 21369 31343 21403
rect 36461 21369 36495 21403
rect 1593 21301 1627 21335
rect 2237 21301 2271 21335
rect 2881 21301 2915 21335
rect 7205 21301 7239 21335
rect 7389 21301 7423 21335
rect 7849 21301 7883 21335
rect 8217 21301 8251 21335
rect 17693 21301 17727 21335
rect 26065 21301 26099 21335
rect 39037 21301 39071 21335
rect 7757 21097 7791 21131
rect 15669 21097 15703 21131
rect 17233 21097 17267 21131
rect 25237 21097 25271 21131
rect 36829 21097 36863 21131
rect 38301 21097 38335 21131
rect 7573 21029 7607 21063
rect 19257 21029 19291 21063
rect 35725 21029 35759 21063
rect 1685 20961 1719 20995
rect 15945 20961 15979 20995
rect 17417 20961 17451 20995
rect 17601 20961 17635 20995
rect 19533 20961 19567 20995
rect 32597 20961 32631 20995
rect 1952 20893 1986 20927
rect 7665 20893 7699 20927
rect 7849 20893 7883 20927
rect 8033 20893 8067 20927
rect 10517 20893 10551 20927
rect 15853 20893 15887 20927
rect 16037 20893 16071 20927
rect 16129 20893 16163 20927
rect 17509 20893 17543 20927
rect 17693 20893 17727 20927
rect 19415 20893 19449 20927
rect 19626 20893 19660 20927
rect 19718 20893 19752 20927
rect 21557 20893 21591 20927
rect 25421 20893 25455 20927
rect 25697 20893 25731 20927
rect 28181 20893 28215 20927
rect 32321 20893 32355 20927
rect 35081 20893 35115 20927
rect 35174 20893 35208 20927
rect 35546 20893 35580 20927
rect 36185 20893 36219 20927
rect 36278 20893 36312 20927
rect 36650 20893 36684 20927
rect 38485 20893 38519 20927
rect 38761 20893 38795 20927
rect 13185 20825 13219 20859
rect 21824 20825 21858 20859
rect 27261 20825 27295 20859
rect 35357 20825 35391 20859
rect 35449 20825 35483 20859
rect 36461 20825 36495 20859
rect 36553 20825 36587 20859
rect 38669 20825 38703 20859
rect 3065 20757 3099 20791
rect 7297 20757 7331 20791
rect 10333 20757 10367 20791
rect 13277 20757 13311 20791
rect 22937 20757 22971 20791
rect 25605 20757 25639 20791
rect 27353 20757 27387 20791
rect 27997 20757 28031 20791
rect 2145 20553 2179 20587
rect 2513 20553 2547 20587
rect 7205 20553 7239 20587
rect 10241 20553 10275 20587
rect 10609 20553 10643 20587
rect 17969 20553 18003 20587
rect 22385 20553 22419 20587
rect 25789 20553 25823 20587
rect 27537 20553 27571 20587
rect 12449 20485 12483 20519
rect 12909 20485 12943 20519
rect 13093 20485 13127 20519
rect 22017 20485 22051 20519
rect 28242 20485 28276 20519
rect 36001 20485 36035 20519
rect 36093 20485 36127 20519
rect 1409 20417 1443 20451
rect 3801 20417 3835 20451
rect 6837 20417 6871 20451
rect 7021 20417 7055 20451
rect 7665 20417 7699 20451
rect 7941 20417 7975 20451
rect 12265 20417 12299 20451
rect 15577 20417 15611 20451
rect 16681 20417 16715 20451
rect 19809 20417 19843 20451
rect 22201 20417 22235 20451
rect 22477 20417 22511 20451
rect 25697 20417 25731 20451
rect 27169 20417 27203 20451
rect 27353 20417 27387 20451
rect 35725 20417 35759 20451
rect 35873 20417 35907 20451
rect 36190 20417 36224 20451
rect 39385 20417 39419 20451
rect 2605 20349 2639 20383
rect 2697 20349 2731 20383
rect 7757 20349 7791 20383
rect 10701 20349 10735 20383
rect 10793 20349 10827 20383
rect 15301 20349 15335 20383
rect 16957 20349 16991 20383
rect 18153 20349 18187 20383
rect 18245 20349 18279 20383
rect 18337 20349 18371 20383
rect 18429 20349 18463 20383
rect 19533 20349 19567 20383
rect 19718 20349 19752 20383
rect 19901 20349 19935 20383
rect 19993 20349 20027 20383
rect 27997 20349 28031 20383
rect 39129 20349 39163 20383
rect 36369 20281 36403 20315
rect 1593 20213 1627 20247
rect 3617 20213 3651 20247
rect 7665 20213 7699 20247
rect 8125 20213 8159 20247
rect 13093 20213 13127 20247
rect 13277 20213 13311 20247
rect 29377 20213 29411 20247
rect 40509 20213 40543 20247
rect 2513 20009 2547 20043
rect 7389 20009 7423 20043
rect 11805 20009 11839 20043
rect 12817 20009 12851 20043
rect 14657 20009 14691 20043
rect 28641 20009 28675 20043
rect 38761 20009 38795 20043
rect 38301 19941 38335 19975
rect 3801 19873 3835 19907
rect 7297 19873 7331 19907
rect 8401 19873 8435 19907
rect 10425 19873 10459 19907
rect 13553 19873 13587 19907
rect 15577 19873 15611 19907
rect 19717 19873 19751 19907
rect 19993 19873 20027 19907
rect 20177 19873 20211 19907
rect 29653 19873 29687 19907
rect 29837 19873 29871 19907
rect 31217 19873 31251 19907
rect 38945 19873 38979 19907
rect 39129 19873 39163 19907
rect 39221 19873 39255 19907
rect 2697 19805 2731 19839
rect 4057 19805 4091 19839
rect 7389 19805 7423 19839
rect 10692 19805 10726 19839
rect 13093 19805 13127 19839
rect 15485 19805 15519 19839
rect 15669 19805 15703 19839
rect 15761 19805 15795 19839
rect 17417 19805 17451 19839
rect 17693 19805 17727 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 24409 19805 24443 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 29561 19805 29595 19839
rect 30757 19805 30791 19839
rect 35817 19805 35851 19839
rect 35965 19805 35999 19839
rect 36282 19805 36316 19839
rect 38025 19805 38059 19839
rect 38301 19805 38335 19839
rect 39037 19805 39071 19839
rect 1869 19737 1903 19771
rect 2053 19737 2087 19771
rect 6929 19737 6963 19771
rect 8033 19737 8067 19771
rect 8217 19737 8251 19771
rect 13001 19737 13035 19771
rect 14473 19737 14507 19771
rect 14673 19737 14707 19771
rect 24676 19737 24710 19771
rect 27261 19737 27295 19771
rect 29837 19737 29871 19771
rect 31462 19737 31496 19771
rect 36093 19737 36127 19771
rect 36185 19737 36219 19771
rect 38209 19737 38243 19771
rect 5181 19669 5215 19703
rect 7573 19669 7607 19703
rect 14841 19669 14875 19703
rect 15301 19669 15335 19703
rect 25789 19669 25823 19703
rect 27353 19669 27387 19703
rect 30573 19669 30607 19703
rect 32597 19669 32631 19703
rect 36461 19669 36495 19703
rect 2053 19465 2087 19499
rect 3801 19465 3835 19499
rect 7205 19465 7239 19499
rect 8125 19465 8159 19499
rect 12817 19465 12851 19499
rect 15117 19465 15151 19499
rect 19441 19465 19475 19499
rect 24685 19465 24719 19499
rect 25053 19465 25087 19499
rect 27353 19465 27387 19499
rect 30573 19465 30607 19499
rect 34069 19465 34103 19499
rect 38761 19465 38795 19499
rect 3709 19397 3743 19431
rect 7665 19397 7699 19431
rect 20545 19397 20579 19431
rect 26065 19397 26099 19431
rect 26265 19397 26299 19431
rect 26985 19397 27019 19431
rect 27185 19397 27219 19431
rect 31309 19397 31343 19431
rect 33793 19397 33827 19431
rect 1593 19329 1627 19363
rect 2237 19329 2271 19363
rect 6653 19329 6687 19363
rect 7021 19329 7055 19363
rect 7849 19329 7883 19363
rect 7941 19329 7975 19363
rect 11529 19329 11563 19363
rect 11713 19329 11747 19363
rect 12265 19329 12299 19363
rect 13277 19329 13311 19363
rect 13461 19329 13495 19363
rect 13553 19329 13587 19363
rect 15301 19329 15335 19363
rect 15485 19329 15519 19363
rect 17141 19329 17175 19363
rect 18429 19329 18463 19363
rect 19809 19329 19843 19363
rect 21833 19329 21867 19363
rect 22100 19329 22134 19363
rect 24869 19329 24903 19363
rect 25145 19329 25179 19363
rect 29469 19329 29503 19363
rect 29653 19329 29687 19363
rect 30205 19329 30239 19363
rect 30389 19329 30423 19363
rect 31217 19329 31251 19363
rect 31401 19329 31435 19363
rect 32137 19329 32171 19363
rect 33425 19329 33459 19363
rect 33518 19329 33552 19363
rect 33701 19329 33735 19363
rect 33890 19329 33924 19363
rect 35541 19329 35575 19363
rect 38945 19329 38979 19363
rect 39129 19329 39163 19363
rect 39221 19329 39255 19363
rect 3893 19261 3927 19295
rect 14013 19261 14047 19295
rect 15393 19261 15427 19295
rect 15577 19261 15611 19295
rect 18153 19261 18187 19295
rect 19625 19261 19659 19295
rect 19717 19261 19751 19295
rect 19901 19261 19935 19295
rect 31033 19261 31067 19295
rect 31585 19261 31619 19295
rect 32413 19261 32447 19295
rect 35265 19261 35299 19295
rect 3341 19193 3375 19227
rect 25789 19193 25823 19227
rect 1409 19125 1443 19159
rect 7021 19125 7055 19159
rect 7665 19125 7699 19159
rect 17233 19125 17267 19159
rect 20637 19125 20671 19159
rect 23213 19125 23247 19159
rect 26249 19125 26283 19159
rect 26433 19125 26467 19159
rect 27169 19125 27203 19159
rect 27721 19125 27755 19159
rect 29561 19125 29595 19159
rect 3157 18921 3191 18955
rect 7205 18921 7239 18955
rect 10425 18921 10459 18955
rect 19533 18921 19567 18955
rect 20545 18921 20579 18955
rect 22201 18921 22235 18955
rect 28825 18921 28859 18955
rect 29009 18921 29043 18955
rect 29561 18921 29595 18955
rect 11989 18853 12023 18887
rect 25421 18853 25455 18887
rect 32689 18853 32723 18887
rect 39865 18853 39899 18887
rect 7113 18785 7147 18819
rect 17417 18785 17451 18819
rect 17693 18785 17727 18819
rect 19993 18785 20027 18819
rect 20821 18785 20855 18819
rect 34713 18785 34747 18819
rect 34989 18785 35023 18819
rect 1777 18717 1811 18751
rect 6837 18717 6871 18751
rect 7849 18717 7883 18751
rect 8033 18717 8067 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 10333 18717 10367 18751
rect 10517 18717 10551 18751
rect 11805 18717 11839 18751
rect 12541 18717 12575 18751
rect 14105 18717 14139 18751
rect 19717 18717 19751 18751
rect 19809 18717 19843 18751
rect 19901 18717 19935 18751
rect 20729 18717 20763 18751
rect 20913 18717 20947 18751
rect 21005 18717 21039 18751
rect 22385 18717 22419 18751
rect 22661 18717 22695 18751
rect 29817 18717 29851 18751
rect 29926 18714 29960 18748
rect 30026 18717 30060 18751
rect 30205 18717 30239 18751
rect 32045 18717 32079 18751
rect 32193 18717 32227 18751
rect 32321 18717 32355 18751
rect 32551 18717 32585 18751
rect 36001 18717 36035 18751
rect 36149 18717 36183 18751
rect 36507 18717 36541 18751
rect 37197 18717 37231 18751
rect 37345 18717 37379 18751
rect 37662 18717 37696 18751
rect 40049 18717 40083 18751
rect 2044 18649 2078 18683
rect 8217 18649 8251 18683
rect 9045 18649 9079 18683
rect 15577 18649 15611 18683
rect 25237 18649 25271 18683
rect 28641 18649 28675 18683
rect 32413 18649 32447 18683
rect 36277 18649 36311 18683
rect 36369 18649 36403 18683
rect 37473 18649 37507 18683
rect 37565 18649 37599 18683
rect 40141 18649 40175 18683
rect 7389 18581 7423 18615
rect 12725 18581 12759 18615
rect 14289 18581 14323 18615
rect 15853 18581 15887 18615
rect 22569 18581 22603 18615
rect 28851 18581 28885 18615
rect 36645 18581 36679 18615
rect 37841 18581 37875 18615
rect 40233 18581 40267 18615
rect 40417 18581 40451 18615
rect 1593 18377 1627 18411
rect 2605 18377 2639 18411
rect 3893 18377 3927 18411
rect 9689 18377 9723 18411
rect 11897 18377 11931 18411
rect 19993 18377 20027 18411
rect 2697 18309 2731 18343
rect 31217 18309 31251 18343
rect 31309 18309 31343 18343
rect 38853 18309 38887 18343
rect 1409 18241 1443 18275
rect 3801 18241 3835 18275
rect 6929 18241 6963 18275
rect 8309 18241 8343 18275
rect 8576 18241 8610 18275
rect 11713 18241 11747 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 17233 18241 17267 18275
rect 18245 18241 18279 18275
rect 18337 18241 18371 18275
rect 19165 18241 19199 18275
rect 19442 18241 19476 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 27077 18241 27111 18275
rect 27333 18241 27367 18275
rect 29009 18241 29043 18275
rect 29193 18241 29227 18275
rect 29285 18241 29319 18275
rect 30941 18241 30975 18275
rect 31089 18241 31123 18275
rect 31447 18241 31481 18275
rect 33609 18241 33643 18275
rect 35173 18241 35207 18275
rect 37289 18241 37323 18275
rect 37473 18241 37507 18275
rect 39681 18241 39715 18275
rect 40765 18241 40799 18275
rect 2881 18173 2915 18207
rect 11529 18173 11563 18207
rect 16865 18173 16899 18207
rect 17049 18173 17083 18207
rect 17141 18173 17175 18207
rect 17325 18173 17359 18207
rect 18061 18173 18095 18207
rect 18153 18173 18187 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 20269 18173 20303 18207
rect 20453 18173 20487 18207
rect 32321 18173 32355 18207
rect 32597 18173 32631 18207
rect 33885 18173 33919 18207
rect 34897 18173 34931 18207
rect 39037 18173 39071 18207
rect 39773 18173 39807 18207
rect 40509 18173 40543 18207
rect 17877 18105 17911 18139
rect 28457 18105 28491 18139
rect 2237 18037 2271 18071
rect 7113 18037 7147 18071
rect 18981 18037 19015 18071
rect 29009 18037 29043 18071
rect 31585 18037 31619 18071
rect 37381 18037 37415 18071
rect 40049 18037 40083 18071
rect 41889 18037 41923 18071
rect 6193 17833 6227 17867
rect 8953 17833 8987 17867
rect 13277 17833 13311 17867
rect 15945 17833 15979 17867
rect 18153 17833 18187 17867
rect 27169 17833 27203 17867
rect 29561 17833 29595 17867
rect 39865 17833 39899 17867
rect 48329 17833 48363 17867
rect 2145 17765 2179 17799
rect 3801 17765 3835 17799
rect 29929 17765 29963 17799
rect 18521 17697 18555 17731
rect 19257 17697 19291 17731
rect 24409 17697 24443 17731
rect 27261 17697 27295 17731
rect 32321 17697 32355 17731
rect 42625 17697 42659 17731
rect 45477 17697 45511 17731
rect 1869 17629 1903 17663
rect 2697 17629 2731 17663
rect 3985 17629 4019 17663
rect 4813 17629 4847 17663
rect 6837 17629 6871 17663
rect 7113 17629 7147 17663
rect 9137 17629 9171 17663
rect 9397 17639 9431 17673
rect 12173 17629 12207 17663
rect 12817 17629 12851 17663
rect 13093 17629 13127 17663
rect 14565 17629 14599 17663
rect 18337 17629 18371 17663
rect 18429 17629 18463 17663
rect 18613 17629 18647 17663
rect 19533 17629 19567 17663
rect 21649 17629 21683 17663
rect 26985 17629 27019 17663
rect 27077 17629 27111 17663
rect 29561 17629 29595 17663
rect 29745 17629 29779 17663
rect 32045 17629 32079 17663
rect 34713 17629 34747 17663
rect 37197 17629 37231 17663
rect 37289 17629 37323 17663
rect 37381 17629 37415 17663
rect 37565 17629 37599 17663
rect 40049 17629 40083 17663
rect 40325 17629 40359 17663
rect 5080 17561 5114 17595
rect 6653 17561 6687 17595
rect 9321 17561 9355 17595
rect 13001 17561 13035 17595
rect 14832 17561 14866 17595
rect 21916 17561 21950 17595
rect 24676 17561 24710 17595
rect 42892 17561 42926 17595
rect 45722 17561 45756 17595
rect 48237 17561 48271 17595
rect 2881 17493 2915 17527
rect 7021 17493 7055 17527
rect 12265 17493 12299 17527
rect 23029 17493 23063 17527
rect 25789 17493 25823 17527
rect 34897 17493 34931 17527
rect 36921 17493 36955 17527
rect 40233 17493 40267 17527
rect 44005 17493 44039 17527
rect 46857 17493 46891 17527
rect 15301 17289 15335 17323
rect 15669 17289 15703 17323
rect 22385 17289 22419 17323
rect 24685 17289 24719 17323
rect 26249 17289 26283 17323
rect 31585 17289 31619 17323
rect 38945 17289 38979 17323
rect 42901 17289 42935 17323
rect 45293 17289 45327 17323
rect 13277 17221 13311 17255
rect 13829 17221 13863 17255
rect 27629 17221 27663 17255
rect 31217 17221 31251 17255
rect 32413 17221 32447 17255
rect 32505 17221 32539 17255
rect 1409 17153 1443 17187
rect 2697 17153 2731 17187
rect 3341 17153 3375 17187
rect 7757 17153 7791 17187
rect 8024 17153 8058 17187
rect 12173 17153 12207 17187
rect 12357 17153 12391 17187
rect 13369 17153 13403 17187
rect 14381 17153 14415 17187
rect 15485 17153 15519 17187
rect 15761 17153 15795 17187
rect 18981 17153 19015 17187
rect 22201 17153 22235 17187
rect 22477 17153 22511 17187
rect 24961 17153 24995 17187
rect 26065 17153 26099 17187
rect 26249 17153 26283 17187
rect 27445 17153 27479 17187
rect 30941 17153 30975 17187
rect 31089 17153 31123 17187
rect 31309 17153 31343 17187
rect 31406 17153 31440 17187
rect 32137 17153 32171 17187
rect 32230 17153 32264 17187
rect 32643 17153 32677 17187
rect 37821 17153 37855 17187
rect 43085 17153 43119 17187
rect 45477 17153 45511 17187
rect 17417 17085 17451 17119
rect 17693 17085 17727 17119
rect 18705 17085 18739 17119
rect 22017 17085 22051 17119
rect 24869 17085 24903 17119
rect 25237 17085 25271 17119
rect 25329 17085 25363 17119
rect 37565 17085 37599 17119
rect 12357 17017 12391 17051
rect 32781 17017 32815 17051
rect 1593 16949 1627 16983
rect 2513 16949 2547 16983
rect 3157 16949 3191 16983
rect 9137 16949 9171 16983
rect 13093 16949 13127 16983
rect 14473 16949 14507 16983
rect 8953 16745 8987 16779
rect 12265 16745 12299 16779
rect 14657 16745 14691 16779
rect 35265 16745 35299 16779
rect 35817 16745 35851 16779
rect 42901 16745 42935 16779
rect 43085 16745 43119 16779
rect 45569 16745 45603 16779
rect 13369 16677 13403 16711
rect 10885 16609 10919 16643
rect 18429 16609 18463 16643
rect 36921 16609 36955 16643
rect 37013 16609 37047 16643
rect 37197 16609 37231 16643
rect 40509 16609 40543 16643
rect 43913 16609 43947 16643
rect 44005 16609 44039 16643
rect 45017 16609 45051 16643
rect 1869 16541 1903 16575
rect 2136 16541 2170 16575
rect 3985 16541 4019 16575
rect 9137 16541 9171 16575
rect 9413 16541 9447 16575
rect 18337 16541 18371 16575
rect 18521 16541 18555 16575
rect 18613 16541 18647 16575
rect 25145 16541 25179 16575
rect 30757 16541 30791 16575
rect 30941 16541 30975 16575
rect 33793 16541 33827 16575
rect 33977 16541 34011 16575
rect 37105 16541 37139 16575
rect 41153 16541 41187 16575
rect 43729 16541 43763 16575
rect 43821 16541 43855 16575
rect 45201 16541 45235 16575
rect 46581 16541 46615 16575
rect 46949 16541 46983 16575
rect 48145 16541 48179 16575
rect 8217 16473 8251 16507
rect 11130 16473 11164 16507
rect 13185 16473 13219 16507
rect 14565 16473 14599 16507
rect 29561 16473 29595 16507
rect 29745 16473 29779 16507
rect 35081 16473 35115 16507
rect 35265 16473 35299 16507
rect 40325 16473 40359 16507
rect 42717 16473 42751 16507
rect 46857 16473 46891 16507
rect 47066 16473 47100 16507
rect 3249 16405 3283 16439
rect 3801 16405 3835 16439
rect 8309 16405 8343 16439
rect 9321 16405 9355 16439
rect 18153 16405 18187 16439
rect 25329 16405 25363 16439
rect 29929 16405 29963 16439
rect 30849 16405 30883 16439
rect 33885 16405 33919 16439
rect 35449 16405 35483 16439
rect 36737 16405 36771 16439
rect 40969 16405 41003 16439
rect 42927 16405 42961 16439
rect 43545 16405 43579 16439
rect 45293 16405 45327 16439
rect 45385 16405 45419 16439
rect 47225 16405 47259 16439
rect 47961 16405 47995 16439
rect 2421 16201 2455 16235
rect 2789 16201 2823 16235
rect 7757 16201 7791 16235
rect 10793 16201 10827 16235
rect 18061 16201 18095 16235
rect 19073 16201 19107 16235
rect 25329 16201 25363 16235
rect 28641 16201 28675 16235
rect 30665 16201 30699 16235
rect 32413 16201 32447 16235
rect 33149 16201 33183 16235
rect 44925 16201 44959 16235
rect 46397 16201 46431 16235
rect 49709 16201 49743 16235
rect 20729 16133 20763 16167
rect 20913 16133 20947 16167
rect 29530 16133 29564 16167
rect 32689 16133 32723 16167
rect 34428 16133 34462 16167
rect 40592 16133 40626 16167
rect 48574 16133 48608 16167
rect 1593 16065 1627 16099
rect 2881 16065 2915 16099
rect 6633 16065 6667 16099
rect 10977 16065 11011 16099
rect 13369 16065 13403 16099
rect 14648 16065 14682 16099
rect 17417 16065 17451 16099
rect 17509 16065 17543 16099
rect 18245 16065 18279 16099
rect 18429 16065 18463 16099
rect 18521 16065 18555 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 21833 16065 21867 16099
rect 22089 16065 22123 16099
rect 23949 16065 23983 16099
rect 24216 16065 24250 16099
rect 28825 16065 28859 16099
rect 31125 16065 31159 16099
rect 32321 16065 32355 16099
rect 32505 16065 32539 16099
rect 33425 16065 33459 16099
rect 33609 16065 33643 16099
rect 34161 16065 34195 16099
rect 40325 16065 40359 16099
rect 43913 16065 43947 16099
rect 44097 16065 44131 16099
rect 44557 16065 44591 16099
rect 44741 16065 44775 16099
rect 46213 16065 46247 16099
rect 46397 16065 46431 16099
rect 46857 16065 46891 16099
rect 47041 16065 47075 16099
rect 47593 16065 47627 16099
rect 48329 16065 48363 16099
rect 3065 15997 3099 16031
rect 6377 15997 6411 16031
rect 14381 15997 14415 16031
rect 17049 15997 17083 16031
rect 17233 15997 17267 16031
rect 17325 15997 17359 16031
rect 18338 15997 18372 16031
rect 19349 15997 19383 16031
rect 19533 15997 19567 16031
rect 29285 15997 29319 16031
rect 33333 15997 33367 16031
rect 33517 15997 33551 16031
rect 47685 15997 47719 16031
rect 15761 15929 15795 15963
rect 32137 15929 32171 15963
rect 46857 15929 46891 15963
rect 1869 15861 1903 15895
rect 13461 15861 13495 15895
rect 20361 15861 20395 15895
rect 20913 15861 20947 15895
rect 21097 15861 21131 15895
rect 23213 15861 23247 15895
rect 31217 15861 31251 15895
rect 35541 15861 35575 15895
rect 41705 15861 41739 15895
rect 44005 15861 44039 15895
rect 6285 15657 6319 15691
rect 10517 15657 10551 15691
rect 14933 15657 14967 15691
rect 16129 15657 16163 15691
rect 18153 15657 18187 15691
rect 19257 15657 19291 15691
rect 24593 15657 24627 15691
rect 26525 15657 26559 15691
rect 30297 15657 30331 15691
rect 33609 15657 33643 15691
rect 33701 15657 33735 15691
rect 35081 15657 35115 15691
rect 40601 15657 40635 15691
rect 54769 15657 54803 15691
rect 2237 15589 2271 15623
rect 16313 15589 16347 15623
rect 26709 15589 26743 15623
rect 30205 15589 30239 15623
rect 37657 15589 37691 15623
rect 2789 15521 2823 15555
rect 11069 15521 11103 15555
rect 15301 15521 15335 15555
rect 15393 15521 15427 15555
rect 18429 15521 18463 15555
rect 18613 15521 18647 15555
rect 19441 15521 19475 15555
rect 19625 15521 19659 15555
rect 25973 15521 26007 15555
rect 33793 15521 33827 15555
rect 35725 15521 35759 15555
rect 40233 15521 40267 15555
rect 41797 15521 41831 15555
rect 41981 15521 42015 15555
rect 42165 15521 42199 15555
rect 1409 15453 1443 15487
rect 2605 15453 2639 15487
rect 3985 15453 4019 15487
rect 6469 15453 6503 15487
rect 6653 15453 6687 15487
rect 6745 15453 6779 15487
rect 10885 15453 10919 15487
rect 15117 15453 15151 15487
rect 15209 15453 15243 15487
rect 18337 15453 18371 15487
rect 18521 15453 18555 15487
rect 19533 15453 19567 15487
rect 19717 15453 19751 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 22293 15453 22327 15487
rect 24777 15453 24811 15487
rect 24961 15453 24995 15487
rect 25053 15453 25087 15487
rect 27353 15453 27387 15487
rect 30113 15453 30147 15487
rect 30297 15453 30331 15487
rect 33517 15453 33551 15487
rect 34897 15453 34931 15487
rect 36001 15453 36035 15487
rect 37933 15453 37967 15487
rect 40417 15453 40451 15487
rect 42073 15453 42107 15487
rect 42257 15453 42291 15487
rect 43545 15453 43579 15487
rect 43729 15453 43763 15487
rect 47041 15453 47075 15487
rect 47133 15453 47167 15487
rect 53389 15453 53423 15487
rect 15945 15385 15979 15419
rect 21833 15385 21867 15419
rect 26341 15385 26375 15419
rect 26541 15385 26575 15419
rect 27169 15385 27203 15419
rect 29929 15385 29963 15419
rect 37657 15385 37691 15419
rect 46857 15385 46891 15419
rect 53634 15385 53668 15419
rect 1593 15317 1627 15351
rect 2697 15317 2731 15351
rect 3801 15317 3835 15351
rect 10977 15317 11011 15351
rect 16155 15317 16189 15351
rect 27537 15317 27571 15351
rect 37841 15317 37875 15351
rect 43729 15317 43763 15351
rect 46949 15317 46983 15351
rect 5641 15113 5675 15147
rect 8677 15113 8711 15147
rect 8769 15113 8803 15147
rect 12081 15113 12115 15147
rect 18061 15113 18095 15147
rect 22845 15113 22879 15147
rect 26985 15113 27019 15147
rect 31493 15113 31527 15147
rect 38761 15113 38795 15147
rect 40969 15113 41003 15147
rect 43637 15113 43671 15147
rect 44281 15113 44315 15147
rect 47685 15113 47719 15147
rect 53021 15113 53055 15147
rect 13461 15045 13495 15079
rect 13645 15045 13679 15079
rect 30941 15045 30975 15079
rect 40877 15045 40911 15079
rect 44097 15045 44131 15079
rect 1961 14977 1995 15011
rect 2228 14977 2262 15011
rect 4261 14977 4295 15011
rect 4528 14977 4562 15011
rect 7389 14977 7423 15011
rect 8861 14977 8895 15011
rect 11989 14977 12023 15011
rect 12633 14977 12667 15011
rect 12817 14977 12851 15011
rect 15301 14977 15335 15011
rect 15485 14977 15519 15011
rect 18429 14977 18463 15011
rect 18521 14977 18555 15011
rect 21005 14977 21039 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22569 14977 22603 15011
rect 27215 14977 27249 15011
rect 27334 14977 27368 15011
rect 27450 14977 27484 15011
rect 27629 14977 27663 15011
rect 28273 14977 28307 15011
rect 30757 14977 30791 15011
rect 31401 14977 31435 15011
rect 31585 14977 31619 15011
rect 34437 14977 34471 15011
rect 37381 14977 37415 15011
rect 37637 14977 37671 15011
rect 43269 14977 43303 15011
rect 43453 14977 43487 15011
rect 44373 14977 44407 15011
rect 47593 14977 47627 15011
rect 47777 14977 47811 15011
rect 53205 14977 53239 15011
rect 7205 14909 7239 14943
rect 8125 14909 8159 14943
rect 8309 14909 8343 14943
rect 14657 14909 14691 14943
rect 15209 14909 15243 14943
rect 15393 14909 15427 14943
rect 18245 14909 18279 14943
rect 18337 14909 18371 14943
rect 3341 14773 3375 14807
rect 7573 14773 7607 14807
rect 12633 14773 12667 14807
rect 13645 14773 13679 14807
rect 13829 14773 13863 14807
rect 15025 14773 15059 14807
rect 21189 14773 21223 14807
rect 21833 14773 21867 14807
rect 28089 14773 28123 14807
rect 34621 14773 34655 14807
rect 43269 14773 43303 14807
rect 44097 14773 44131 14807
rect 2697 14569 2731 14603
rect 5181 14569 5215 14603
rect 15761 14569 15795 14603
rect 16405 14569 16439 14603
rect 16589 14569 16623 14603
rect 18153 14569 18187 14603
rect 26709 14569 26743 14603
rect 31953 14569 31987 14603
rect 33701 14569 33735 14603
rect 36185 14569 36219 14603
rect 37381 14569 37415 14603
rect 37473 14569 37507 14603
rect 40141 14569 40175 14603
rect 43637 14569 43671 14603
rect 43729 14501 43763 14535
rect 1409 14433 1443 14467
rect 1685 14433 1719 14467
rect 12265 14433 12299 14467
rect 12725 14433 12759 14467
rect 14381 14433 14415 14467
rect 18429 14433 18463 14467
rect 18521 14433 18555 14467
rect 22017 14433 22051 14467
rect 25237 14433 25271 14467
rect 30757 14433 30791 14467
rect 31033 14433 31067 14467
rect 40325 14433 40359 14467
rect 43913 14433 43947 14467
rect 2881 14365 2915 14399
rect 5365 14365 5399 14399
rect 5641 14365 5675 14399
rect 7481 14365 7515 14399
rect 7573 14365 7607 14399
rect 7757 14365 7791 14399
rect 10517 14365 10551 14399
rect 10793 14365 10827 14399
rect 11161 14365 11195 14399
rect 12817 14365 12851 14399
rect 14648 14365 14682 14399
rect 18337 14365 18371 14399
rect 18613 14365 18647 14399
rect 21649 14365 21683 14399
rect 21741 14365 21775 14399
rect 26617 14365 26651 14399
rect 26801 14365 26835 14399
rect 27261 14365 27295 14399
rect 27528 14365 27562 14399
rect 30849 14365 30883 14399
rect 30941 14365 30975 14399
rect 31585 14365 31619 14399
rect 31769 14365 31803 14399
rect 33517 14365 33551 14399
rect 36093 14365 36127 14399
rect 37013 14365 37047 14399
rect 37105 14365 37139 14399
rect 37473 14365 37507 14399
rect 40049 14365 40083 14399
rect 43637 14365 43671 14399
rect 46581 14365 46615 14399
rect 50169 14365 50203 14399
rect 53665 14365 53699 14399
rect 53849 14365 53883 14399
rect 7665 14297 7699 14331
rect 16221 14297 16255 14331
rect 16437 14297 16471 14331
rect 22109 14297 22143 14331
rect 25053 14297 25087 14331
rect 46826 14297 46860 14331
rect 50436 14297 50470 14331
rect 5549 14229 5583 14263
rect 7941 14229 7975 14263
rect 11805 14229 11839 14263
rect 12449 14229 12483 14263
rect 21465 14229 21499 14263
rect 28641 14229 28675 14263
rect 30573 14229 30607 14263
rect 36553 14229 36587 14263
rect 37197 14229 37231 14263
rect 40601 14229 40635 14263
rect 47961 14229 47995 14263
rect 51549 14229 51583 14263
rect 53757 14229 53791 14263
rect 2145 14025 2179 14059
rect 3249 14025 3283 14059
rect 10977 14025 11011 14059
rect 14795 14025 14829 14059
rect 23213 14025 23247 14059
rect 31585 14025 31619 14059
rect 32321 14025 32355 14059
rect 40233 14025 40267 14059
rect 46673 14025 46707 14059
rect 50629 14025 50663 14059
rect 10609 13957 10643 13991
rect 22078 13957 22112 13991
rect 24654 13957 24688 13991
rect 27997 13957 28031 13991
rect 30450 13957 30484 13991
rect 40141 13957 40175 13991
rect 40969 13957 41003 13991
rect 45477 13957 45511 13991
rect 53472 13957 53506 13991
rect 1409 13889 1443 13923
rect 2329 13889 2363 13923
rect 3157 13889 3191 13923
rect 7849 13889 7883 13923
rect 8217 13889 8251 13923
rect 8401 13889 8435 13923
rect 8953 13889 8987 13923
rect 10793 13889 10827 13923
rect 11989 13889 12023 13923
rect 21833 13889 21867 13923
rect 24409 13889 24443 13923
rect 27813 13889 27847 13923
rect 32137 13889 32171 13923
rect 33701 13889 33735 13923
rect 34069 13889 34103 13923
rect 34796 13889 34830 13923
rect 36553 13889 36587 13923
rect 36737 13889 36771 13923
rect 40785 13889 40819 13923
rect 41061 13889 41095 13923
rect 45293 13889 45327 13923
rect 46581 13889 46615 13923
rect 50537 13889 50571 13923
rect 50721 13889 50755 13923
rect 3341 13821 3375 13855
rect 12265 13821 12299 13855
rect 13277 13821 13311 13855
rect 13553 13821 13587 13855
rect 14565 13821 14599 13855
rect 30205 13821 30239 13855
rect 34529 13821 34563 13855
rect 36645 13821 36679 13855
rect 45109 13821 45143 13855
rect 46857 13821 46891 13855
rect 53205 13821 53239 13855
rect 40785 13753 40819 13787
rect 1593 13685 1627 13719
rect 2789 13685 2823 13719
rect 9045 13685 9079 13719
rect 25789 13685 25823 13719
rect 35909 13685 35943 13719
rect 46213 13685 46247 13719
rect 54585 13685 54619 13719
rect 6929 13481 6963 13515
rect 11069 13481 11103 13515
rect 28181 13481 28215 13515
rect 28825 13481 28859 13515
rect 30481 13481 30515 13515
rect 32321 13481 32355 13515
rect 33425 13481 33459 13515
rect 35081 13481 35115 13515
rect 36369 13481 36403 13515
rect 36645 13481 36679 13515
rect 40233 13481 40267 13515
rect 44097 13481 44131 13515
rect 44465 13481 44499 13515
rect 46213 13481 46247 13515
rect 50445 13481 50479 13515
rect 54585 13481 54619 13515
rect 5181 13413 5215 13447
rect 10333 13413 10367 13447
rect 18705 13413 18739 13447
rect 3801 13345 3835 13379
rect 7389 13345 7423 13379
rect 10057 13345 10091 13379
rect 20545 13345 20579 13379
rect 41153 13345 41187 13379
rect 44189 13345 44223 13379
rect 50537 13345 50571 13379
rect 54493 13345 54527 13379
rect 54677 13345 54711 13379
rect 3065 13277 3099 13311
rect 6561 13277 6595 13311
rect 7665 13277 7699 13311
rect 10977 13277 11011 13311
rect 14105 13277 14139 13311
rect 17325 13277 17359 13311
rect 19809 13277 19843 13311
rect 20269 13277 20303 13311
rect 21281 13277 21315 13311
rect 21557 13277 21591 13311
rect 22569 13277 22603 13311
rect 22753 13277 22787 13311
rect 24593 13277 24627 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 28733 13277 28767 13311
rect 28917 13277 28951 13311
rect 30665 13277 30699 13311
rect 30941 13277 30975 13311
rect 32137 13277 32171 13311
rect 35265 13277 35299 13311
rect 35541 13277 35575 13311
rect 36185 13277 36219 13311
rect 39957 13277 39991 13311
rect 41420 13277 41454 13311
rect 44281 13277 44315 13311
rect 46213 13277 46247 13311
rect 46397 13277 46431 13311
rect 49157 13277 49191 13311
rect 49341 13277 49375 13311
rect 50261 13277 50295 13311
rect 50353 13277 50387 13311
rect 53665 13277 53699 13311
rect 53757 13277 53791 13311
rect 54401 13277 54435 13311
rect 1869 13209 1903 13243
rect 2237 13209 2271 13243
rect 4046 13209 4080 13243
rect 6745 13209 6779 13243
rect 17592 13209 17626 13243
rect 28089 13209 28123 13243
rect 33149 13209 33183 13243
rect 35449 13209 35483 13243
rect 43821 13209 43855 13243
rect 2881 13141 2915 13175
rect 10517 13141 10551 13175
rect 14289 13141 14323 13175
rect 22753 13141 22787 13175
rect 24777 13141 24811 13175
rect 30849 13141 30883 13175
rect 40417 13141 40451 13175
rect 42533 13141 42567 13175
rect 49249 13141 49283 13175
rect 53941 13141 53975 13175
rect 7205 12937 7239 12971
rect 9965 12937 9999 12971
rect 17969 12937 18003 12971
rect 18337 12937 18371 12971
rect 21005 12937 21039 12971
rect 24409 12937 24443 12971
rect 48053 12937 48087 12971
rect 50997 12937 51031 12971
rect 57253 12937 57287 12971
rect 13277 12869 13311 12903
rect 15301 12869 15335 12903
rect 15517 12869 15551 12903
rect 19993 12869 20027 12903
rect 20821 12869 20855 12903
rect 28365 12869 28399 12903
rect 29469 12869 29503 12903
rect 29561 12869 29595 12903
rect 38577 12869 38611 12903
rect 44649 12869 44683 12903
rect 47961 12869 47995 12903
rect 49056 12869 49090 12903
rect 1409 12801 1443 12835
rect 2697 12801 2731 12835
rect 3341 12801 3375 12835
rect 7205 12801 7239 12835
rect 7849 12801 7883 12835
rect 8585 12801 8619 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10517 12801 10551 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 12449 12801 12483 12835
rect 13369 12801 13403 12835
rect 15025 12801 15059 12835
rect 18172 12801 18206 12835
rect 18429 12801 18463 12835
rect 20177 12801 20211 12835
rect 24133 12801 24167 12835
rect 28089 12801 28123 12835
rect 28237 12801 28271 12835
rect 28457 12801 28491 12835
rect 28595 12801 28629 12835
rect 29193 12801 29227 12835
rect 29341 12801 29375 12835
rect 29658 12801 29692 12835
rect 38761 12801 38795 12835
rect 39773 12801 39807 12835
rect 39957 12801 39991 12835
rect 40969 12801 41003 12835
rect 43913 12801 43947 12835
rect 44097 12801 44131 12835
rect 44281 12801 44315 12835
rect 45569 12801 45603 12835
rect 50813 12801 50847 12835
rect 53665 12801 53699 12835
rect 53849 12801 53883 12835
rect 53941 12801 53975 12835
rect 54677 12801 54711 12835
rect 56129 12801 56163 12835
rect 8309 12733 8343 12767
rect 12633 12733 12667 12767
rect 24409 12733 24443 12767
rect 41245 12733 41279 12767
rect 48789 12733 48823 12767
rect 50629 12733 50663 12767
rect 54953 12733 54987 12767
rect 55873 12733 55907 12767
rect 3157 12665 3191 12699
rect 11805 12665 11839 12699
rect 13093 12665 13127 12699
rect 20453 12665 20487 12699
rect 29837 12665 29871 12699
rect 44649 12665 44683 12699
rect 50169 12665 50203 12699
rect 1593 12597 1627 12631
rect 2513 12597 2547 12631
rect 10885 12597 10919 12631
rect 13553 12597 13587 12631
rect 15485 12597 15519 12631
rect 15669 12597 15703 12631
rect 21005 12597 21039 12631
rect 21189 12597 21223 12631
rect 24225 12597 24259 12631
rect 28733 12597 28767 12631
rect 38945 12597 38979 12631
rect 40141 12597 40175 12631
rect 45385 12597 45419 12631
rect 53941 12597 53975 12631
rect 54769 12597 54803 12631
rect 54861 12597 54895 12631
rect 2329 12393 2363 12427
rect 5917 12393 5951 12427
rect 21925 12393 21959 12427
rect 32597 12393 32631 12427
rect 39221 12393 39255 12427
rect 46673 12393 46707 12427
rect 48973 12393 49007 12427
rect 50445 12393 50479 12427
rect 50629 12393 50663 12427
rect 55321 12393 55355 12427
rect 10057 12325 10091 12359
rect 11069 12325 11103 12359
rect 22753 12325 22787 12359
rect 26617 12325 26651 12359
rect 33333 12325 33367 12359
rect 40049 12325 40083 12359
rect 43637 12325 43671 12359
rect 2881 12257 2915 12291
rect 4445 12257 4479 12291
rect 9321 12257 9355 12291
rect 9413 12257 9447 12291
rect 22017 12257 22051 12291
rect 27721 12257 27755 12291
rect 28089 12257 28123 12291
rect 35909 12257 35943 12291
rect 45293 12257 45327 12291
rect 49065 12257 49099 12291
rect 51457 12257 51491 12291
rect 53941 12257 53975 12291
rect 1593 12189 1627 12223
rect 4261 12189 4295 12223
rect 6193 12189 6227 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 9137 12189 9171 12223
rect 9873 12189 9907 12223
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 14473 12189 14507 12223
rect 17877 12189 17911 12223
rect 18153 12189 18187 12223
rect 21925 12189 21959 12223
rect 22937 12189 22971 12223
rect 23029 12189 23063 12223
rect 25973 12189 26007 12223
rect 26066 12189 26100 12223
rect 26249 12189 26283 12223
rect 26438 12189 26472 12223
rect 28365 12189 28399 12223
rect 31585 12189 31619 12223
rect 32321 12189 32355 12223
rect 32413 12189 32447 12223
rect 33333 12189 33367 12223
rect 35817 12189 35851 12223
rect 36645 12189 36679 12223
rect 36737 12189 36771 12223
rect 36921 12189 36955 12223
rect 37013 12189 37047 12223
rect 37657 12189 37691 12223
rect 37841 12189 37875 12223
rect 37933 12189 37967 12223
rect 39129 12189 39163 12223
rect 39313 12189 39347 12223
rect 39871 12189 39905 12223
rect 40693 12189 40727 12223
rect 45560 12189 45594 12223
rect 48789 12189 48823 12223
rect 48881 12189 48915 12223
rect 51641 12189 51675 12223
rect 53757 12189 53791 12223
rect 53849 12189 53883 12223
rect 54033 12189 54067 12223
rect 55597 12189 55631 12223
rect 2789 12121 2823 12155
rect 5549 12121 5583 12155
rect 8217 12121 8251 12155
rect 8401 12121 8435 12155
rect 14740 12121 14774 12155
rect 22753 12121 22787 12155
rect 26341 12121 26375 12155
rect 31769 12121 31803 12155
rect 43269 12121 43303 12155
rect 44281 12121 44315 12155
rect 50261 12121 50295 12155
rect 51733 12121 51767 12155
rect 55321 12121 55355 12155
rect 55505 12121 55539 12155
rect 1409 12053 1443 12087
rect 2697 12053 2731 12087
rect 5926 12053 5960 12087
rect 7205 12053 7239 12087
rect 8953 12053 8987 12087
rect 15853 12053 15887 12087
rect 22293 12053 22327 12087
rect 36461 12053 36495 12087
rect 37473 12053 37507 12087
rect 40785 12053 40819 12087
rect 43729 12053 43763 12087
rect 44373 12053 44407 12087
rect 50471 12053 50505 12087
rect 51825 12053 51859 12087
rect 52009 12053 52043 12087
rect 53573 12053 53607 12087
rect 3985 11849 4019 11883
rect 7205 11849 7239 11883
rect 8861 11849 8895 11883
rect 15117 11849 15151 11883
rect 21103 11849 21137 11883
rect 25973 11849 26007 11883
rect 27353 11849 27387 11883
rect 27537 11849 27571 11883
rect 53389 11849 53423 11883
rect 53957 11849 53991 11883
rect 54125 11849 54159 11883
rect 55229 11849 55263 11883
rect 11897 11781 11931 11815
rect 13737 11781 13771 11815
rect 22100 11781 22134 11815
rect 25605 11781 25639 11815
rect 29929 11781 29963 11815
rect 33977 11781 34011 11815
rect 34193 11781 34227 11815
rect 37289 11781 37323 11815
rect 37505 11781 37539 11815
rect 44741 11781 44775 11815
rect 44957 11781 44991 11815
rect 48513 11781 48547 11815
rect 51457 11781 51491 11815
rect 51657 11781 51691 11815
rect 53757 11781 53791 11815
rect 56118 11781 56152 11815
rect 1593 11713 1627 11747
rect 2605 11713 2639 11747
rect 2872 11713 2906 11747
rect 7021 11713 7055 11747
rect 7389 11713 7423 11747
rect 7573 11713 7607 11747
rect 8217 11713 8251 11747
rect 8677 11713 8711 11747
rect 10149 11713 10183 11747
rect 10333 11713 10367 11747
rect 11529 11713 11563 11747
rect 11622 11713 11656 11747
rect 11805 11713 11839 11747
rect 11994 11713 12028 11747
rect 13645 11713 13679 11747
rect 15301 11713 15335 11747
rect 15577 11713 15611 11747
rect 17601 11713 17635 11747
rect 18521 11713 18555 11747
rect 21005 11713 21039 11747
rect 21189 11713 21223 11747
rect 21281 11713 21315 11747
rect 21833 11713 21867 11747
rect 25329 11713 25363 11747
rect 25477 11713 25511 11747
rect 25697 11713 25731 11747
rect 25794 11713 25828 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 27261 11713 27295 11747
rect 32137 11713 32171 11747
rect 34805 11713 34839 11747
rect 35072 11713 35106 11747
rect 38301 11713 38335 11747
rect 38577 11713 38611 11747
rect 39221 11713 39255 11747
rect 39313 11713 39347 11747
rect 40233 11713 40267 11747
rect 40325 11713 40359 11747
rect 40601 11713 40635 11747
rect 41383 11713 41417 11747
rect 41518 11713 41552 11747
rect 41613 11713 41647 11747
rect 41809 11713 41843 11747
rect 42697 11713 42731 11747
rect 48145 11713 48179 11747
rect 55413 11713 55447 11747
rect 55873 11713 55907 11747
rect 8585 11645 8619 11679
rect 10241 11645 10275 11679
rect 13829 11645 13863 11679
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 17417 11645 17451 11679
rect 17509 11645 17543 11679
rect 17693 11645 17727 11679
rect 18245 11645 18279 11679
rect 28549 11645 28583 11679
rect 28825 11645 28859 11679
rect 32413 11645 32447 11679
rect 40509 11645 40543 11679
rect 41153 11645 41187 11679
rect 42441 11645 42475 11679
rect 17233 11577 17267 11611
rect 23213 11577 23247 11611
rect 36185 11577 36219 11611
rect 39497 11577 39531 11611
rect 40693 11577 40727 11611
rect 43821 11577 43855 11611
rect 45109 11577 45143 11611
rect 1409 11509 1443 11543
rect 7389 11509 7423 11543
rect 8677 11509 8711 11543
rect 12173 11509 12207 11543
rect 13277 11509 13311 11543
rect 30205 11509 30239 11543
rect 32229 11509 32263 11543
rect 32321 11509 32355 11543
rect 34161 11509 34195 11543
rect 34345 11509 34379 11543
rect 37473 11509 37507 11543
rect 37657 11509 37691 11543
rect 38393 11509 38427 11543
rect 44925 11509 44959 11543
rect 48513 11509 48547 11543
rect 48697 11509 48731 11543
rect 51641 11509 51675 11543
rect 51825 11509 51859 11543
rect 53941 11509 53975 11543
rect 57253 11509 57287 11543
rect 10609 11305 10643 11339
rect 12357 11305 12391 11339
rect 16221 11305 16255 11339
rect 18061 11305 18095 11339
rect 22385 11305 22419 11339
rect 22569 11305 22603 11339
rect 23857 11305 23891 11339
rect 27721 11305 27755 11339
rect 32505 11305 32539 11339
rect 33333 11305 33367 11339
rect 35173 11305 35207 11339
rect 35541 11305 35575 11339
rect 50905 11305 50939 11339
rect 51089 11305 51123 11339
rect 1593 11237 1627 11271
rect 11621 11237 11655 11271
rect 16405 11237 16439 11271
rect 25421 11237 25455 11271
rect 33425 11237 33459 11271
rect 6469 11169 6503 11203
rect 15209 11169 15243 11203
rect 15485 11169 15519 11203
rect 18245 11169 18279 11203
rect 18337 11169 18371 11203
rect 18521 11169 18555 11203
rect 31125 11169 31159 11203
rect 35633 11169 35667 11203
rect 40969 11169 41003 11203
rect 1409 11101 1443 11135
rect 2421 11101 2455 11135
rect 3065 11101 3099 11135
rect 6101 11101 6135 11135
rect 6377 11101 6411 11135
rect 6653 11101 6687 11135
rect 7113 11101 7147 11135
rect 7389 11101 7423 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 12173 11101 12207 11135
rect 15301 11101 15335 11135
rect 15393 11101 15427 11135
rect 18429 11101 18463 11135
rect 19257 11101 19291 11135
rect 23213 11101 23247 11135
rect 23361 11101 23395 11135
rect 23719 11101 23753 11135
rect 24501 11101 24535 11135
rect 24593 11101 24627 11135
rect 24777 11101 24811 11135
rect 25605 11101 25639 11135
rect 26341 11101 26375 11135
rect 26597 11101 26631 11135
rect 31392 11101 31426 11135
rect 32965 11101 32999 11135
rect 33425 11101 33459 11135
rect 35357 11101 35391 11135
rect 36277 11101 36311 11135
rect 36369 11101 36403 11135
rect 36553 11101 36587 11135
rect 36645 11101 36679 11135
rect 41153 11101 41187 11135
rect 47777 11117 47811 11151
rect 48237 11101 48271 11135
rect 48493 11101 48527 11135
rect 53481 11101 53515 11135
rect 10977 11033 11011 11067
rect 11621 11033 11655 11067
rect 16037 11033 16071 11067
rect 16237 11033 16271 11067
rect 19524 11033 19558 11067
rect 22201 11033 22235 11067
rect 22417 11033 22451 11067
rect 23489 11033 23523 11067
rect 23581 11033 23615 11067
rect 41337 11033 41371 11067
rect 50721 11033 50755 11067
rect 2237 10965 2271 10999
rect 2881 10965 2915 10999
rect 12081 10965 12115 10999
rect 15025 10965 15059 10999
rect 20637 10965 20671 10999
rect 33057 10965 33091 10999
rect 33149 10965 33183 10999
rect 36093 10965 36127 10999
rect 47593 10965 47627 10999
rect 49617 10965 49651 10999
rect 50921 10965 50955 10999
rect 53573 10965 53607 10999
rect 6929 10761 6963 10795
rect 31493 10761 31527 10795
rect 48881 10761 48915 10795
rect 50261 10761 50295 10795
rect 54401 10761 54435 10795
rect 12081 10693 12115 10727
rect 14556 10693 14590 10727
rect 17325 10693 17359 10727
rect 19165 10693 19199 10727
rect 19533 10693 19567 10727
rect 49893 10693 49927 10727
rect 50093 10693 50127 10727
rect 1593 10625 1627 10659
rect 2053 10625 2087 10659
rect 2320 10625 2354 10659
rect 7113 10625 7147 10659
rect 7389 10625 7423 10659
rect 7573 10625 7607 10659
rect 8125 10625 8159 10659
rect 11621 10625 11655 10659
rect 11805 10625 11839 10659
rect 12357 10625 12391 10659
rect 14289 10625 14323 10659
rect 17141 10625 17175 10659
rect 19349 10625 19383 10659
rect 19625 10625 19659 10659
rect 30941 10625 30975 10659
rect 31309 10625 31343 10659
rect 36093 10625 36127 10659
rect 36369 10625 36403 10659
rect 36553 10625 36587 10659
rect 42901 10625 42935 10659
rect 49249 10625 49283 10659
rect 49341 10625 49375 10659
rect 53288 10625 53322 10659
rect 7297 10557 7331 10591
rect 8309 10557 8343 10591
rect 49065 10557 49099 10591
rect 49157 10557 49191 10591
rect 53021 10557 53055 10591
rect 7205 10489 7239 10523
rect 1409 10421 1443 10455
rect 3433 10421 3467 10455
rect 15669 10421 15703 10455
rect 31309 10421 31343 10455
rect 35909 10421 35943 10455
rect 42717 10421 42751 10455
rect 50077 10421 50111 10455
rect 2237 10217 2271 10251
rect 6193 10217 6227 10251
rect 15025 10217 15059 10251
rect 18153 10217 18187 10251
rect 34897 10217 34931 10251
rect 36093 10217 36127 10251
rect 42349 10217 42383 10251
rect 47685 10217 47719 10251
rect 53297 10217 53331 10251
rect 12081 10149 12115 10183
rect 15209 10149 15243 10183
rect 2789 10081 2823 10115
rect 4813 10081 4847 10115
rect 7113 10081 7147 10115
rect 42993 10081 43027 10115
rect 45661 10081 45695 10115
rect 53297 10081 53331 10115
rect 2605 10013 2639 10047
rect 6929 10013 6963 10047
rect 7205 10013 7239 10047
rect 11437 10013 11471 10047
rect 11585 10013 11619 10047
rect 11713 10013 11747 10047
rect 11902 10013 11936 10047
rect 17325 10013 17359 10047
rect 26065 10013 26099 10047
rect 26341 10013 26375 10047
rect 32137 10013 32171 10047
rect 32413 10013 32447 10047
rect 32505 10013 32539 10047
rect 34713 10013 34747 10047
rect 35725 10013 35759 10047
rect 38577 10013 38611 10047
rect 40969 10013 41003 10047
rect 41245 10013 41279 10047
rect 41337 10013 41371 10047
rect 41981 10013 42015 10047
rect 42165 10013 42199 10047
rect 43249 10013 43283 10047
rect 47593 10013 47627 10047
rect 53113 10013 53147 10047
rect 53205 10013 53239 10047
rect 5080 9945 5114 9979
rect 11805 9945 11839 9979
rect 14841 9945 14875 9979
rect 15057 9945 15091 9979
rect 18061 9945 18095 9979
rect 32321 9945 32355 9979
rect 36093 9945 36127 9979
rect 41153 9945 41187 9979
rect 45906 9945 45940 9979
rect 52929 9945 52963 9979
rect 2697 9877 2731 9911
rect 6745 9877 6779 9911
rect 17417 9877 17451 9911
rect 25881 9877 25915 9911
rect 26249 9877 26283 9911
rect 32689 9877 32723 9911
rect 36277 9877 36311 9911
rect 38393 9877 38427 9911
rect 41521 9877 41555 9911
rect 44373 9877 44407 9911
rect 47041 9877 47075 9911
rect 6745 9673 6779 9707
rect 41521 9673 41555 9707
rect 50721 9673 50755 9707
rect 56333 9673 56367 9707
rect 6377 9605 6411 9639
rect 8125 9605 8159 9639
rect 11989 9605 12023 9639
rect 12173 9605 12207 9639
rect 25228 9605 25262 9639
rect 28448 9605 28482 9639
rect 33333 9605 33367 9639
rect 38117 9605 38151 9639
rect 39313 9605 39347 9639
rect 41245 9605 41279 9639
rect 45477 9605 45511 9639
rect 45661 9605 45695 9639
rect 50261 9605 50295 9639
rect 53389 9605 53423 9639
rect 1409 9537 1443 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 9873 9537 9907 9571
rect 13277 9537 13311 9571
rect 13369 9537 13403 9571
rect 14289 9537 14323 9571
rect 16681 9537 16715 9571
rect 18245 9537 18279 9571
rect 19257 9537 19291 9571
rect 19524 9537 19558 9571
rect 22376 9537 22410 9571
rect 30021 9537 30055 9571
rect 31401 9537 31435 9571
rect 33149 9537 33183 9571
rect 33425 9537 33459 9571
rect 33517 9537 33551 9571
rect 34331 9535 34365 9569
rect 35541 9537 35575 9571
rect 35725 9537 35759 9571
rect 37953 9537 37987 9571
rect 38201 9537 38235 9571
rect 38347 9537 38381 9571
rect 39129 9537 39163 9571
rect 40969 9537 41003 9571
rect 41153 9537 41187 9571
rect 41337 9537 41371 9571
rect 42625 9537 42659 9571
rect 45753 9537 45787 9571
rect 48697 9537 48731 9571
rect 48881 9537 48915 9571
rect 49341 9537 49375 9571
rect 50905 9537 50939 9571
rect 51549 9537 51583 9571
rect 52745 9537 52779 9571
rect 52929 9537 52963 9571
rect 53573 9537 53607 9571
rect 54493 9537 54527 9571
rect 55209 9537 55243 9571
rect 13093 9469 13127 9503
rect 14565 9469 14599 9503
rect 16957 9469 16991 9503
rect 18153 9469 18187 9503
rect 18337 9469 18371 9503
rect 18429 9469 18463 9503
rect 22109 9469 22143 9503
rect 24961 9469 24995 9503
rect 28181 9469 28215 9503
rect 31217 9469 31251 9503
rect 34161 9469 34195 9503
rect 38945 9469 38979 9503
rect 42441 9469 42475 9503
rect 48513 9469 48547 9503
rect 49525 9469 49559 9503
rect 50445 9469 50479 9503
rect 50537 9469 50571 9503
rect 50813 9469 50847 9503
rect 51365 9469 51399 9503
rect 51733 9469 51767 9503
rect 54953 9469 54987 9503
rect 26341 9401 26375 9435
rect 33701 9401 33735 9435
rect 38485 9401 38519 9435
rect 45477 9401 45511 9435
rect 54309 9401 54343 9435
rect 1593 9333 1627 9367
rect 8217 9333 8251 9367
rect 8861 9333 8895 9367
rect 9689 9333 9723 9367
rect 13553 9333 13587 9367
rect 17969 9333 18003 9367
rect 20637 9333 20671 9367
rect 23489 9333 23523 9367
rect 29561 9333 29595 9367
rect 30205 9333 30239 9367
rect 31585 9333 31619 9367
rect 32873 9333 32907 9367
rect 34529 9333 34563 9367
rect 35909 9333 35943 9367
rect 42809 9333 42843 9367
rect 52837 9333 52871 9367
rect 53757 9333 53791 9367
rect 2697 9129 2731 9163
rect 10977 9129 11011 9163
rect 17601 9129 17635 9163
rect 20085 9129 20119 9163
rect 22569 9129 22603 9163
rect 25881 9129 25915 9163
rect 31861 9129 31895 9163
rect 35449 9129 35483 9163
rect 41797 9129 41831 9163
rect 52285 9129 52319 9163
rect 53849 9129 53883 9163
rect 54033 9129 54067 9163
rect 36369 9061 36403 9095
rect 50169 9061 50203 9095
rect 1685 8993 1719 9027
rect 14289 8993 14323 9027
rect 16957 8993 16991 9027
rect 17049 8993 17083 9027
rect 17785 8993 17819 9027
rect 17969 8993 18003 9027
rect 18061 8993 18095 9027
rect 20269 8993 20303 9027
rect 20637 8993 20671 9027
rect 21281 8993 21315 9027
rect 22753 8993 22787 9027
rect 23765 8993 23799 9027
rect 25605 8993 25639 9027
rect 32505 8993 32539 9027
rect 42441 8993 42475 9027
rect 1409 8925 1443 8959
rect 2881 8925 2915 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 7205 8925 7239 8959
rect 7481 8925 7515 8959
rect 9597 8925 9631 8959
rect 9853 8925 9887 8959
rect 12357 8925 12391 8959
rect 12541 8925 12575 8959
rect 14381 8925 14415 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17877 8925 17911 8959
rect 20361 8925 20395 8959
rect 21189 8925 21223 8959
rect 21373 8925 21407 8959
rect 22845 8925 22879 8959
rect 23673 8925 23707 8959
rect 23857 8925 23891 8959
rect 25513 8925 25547 8959
rect 30021 8925 30055 8959
rect 34161 8925 34195 8959
rect 35357 8925 35391 8959
rect 37933 8925 37967 8959
rect 38189 8925 38223 8959
rect 45201 8925 45235 8959
rect 50353 8925 50387 8959
rect 50445 8925 50479 8959
rect 52193 8925 52227 8959
rect 20729 8857 20763 8891
rect 23121 8857 23155 8891
rect 23213 8857 23247 8891
rect 30288 8857 30322 8891
rect 32229 8857 32263 8891
rect 36093 8857 36127 8891
rect 50169 8857 50203 8891
rect 53665 8857 53699 8891
rect 53865 8857 53899 8891
rect 3801 8789 3835 8823
rect 4169 8789 4203 8823
rect 7021 8789 7055 8823
rect 7389 8789 7423 8823
rect 14105 8789 14139 8823
rect 16589 8789 16623 8823
rect 31401 8789 31435 8823
rect 32321 8789 32355 8823
rect 33977 8789 34011 8823
rect 39313 8789 39347 8823
rect 42165 8789 42199 8823
rect 42257 8789 42291 8823
rect 45017 8789 45051 8823
rect 2053 8585 2087 8619
rect 7757 8585 7791 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 16681 8585 16715 8619
rect 30941 8585 30975 8619
rect 38577 8585 38611 8619
rect 39037 8585 39071 8619
rect 42441 8585 42475 8619
rect 50721 8585 50755 8619
rect 1777 8517 1811 8551
rect 2872 8517 2906 8551
rect 6644 8517 6678 8551
rect 28089 8517 28123 8551
rect 28305 8517 28339 8551
rect 34130 8517 34164 8551
rect 40325 8517 40359 8551
rect 45722 8517 45756 8551
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 13737 8449 13771 8483
rect 14473 8449 14507 8483
rect 15761 8449 15795 8483
rect 15853 8449 15887 8483
rect 16957 8449 16991 8483
rect 23581 8449 23615 8483
rect 23673 8449 23707 8483
rect 27445 8449 27479 8483
rect 27629 8449 27663 8483
rect 31125 8449 31159 8483
rect 36093 8449 36127 8483
rect 37473 8449 37507 8483
rect 38945 8449 38979 8483
rect 40141 8449 40175 8483
rect 40233 8449 40267 8483
rect 40463 8449 40497 8483
rect 42809 8449 42843 8483
rect 45477 8449 45511 8483
rect 49341 8449 49375 8483
rect 49608 8449 49642 8483
rect 53113 8449 53147 8483
rect 2605 8381 2639 8415
rect 6377 8381 6411 8415
rect 10149 8381 10183 8415
rect 10333 8381 10367 8415
rect 14381 8381 14415 8415
rect 14565 8381 14599 8415
rect 14657 8381 14691 8415
rect 15945 8381 15979 8415
rect 16037 8381 16071 8415
rect 16865 8381 16899 8415
rect 17049 8381 17083 8415
rect 17141 8381 17175 8415
rect 23857 8381 23891 8415
rect 33885 8381 33919 8415
rect 39129 8381 39163 8415
rect 40601 8381 40635 8415
rect 42901 8381 42935 8415
rect 42993 8381 43027 8415
rect 53021 8381 53055 8415
rect 3985 8313 4019 8347
rect 13001 8313 13035 8347
rect 14197 8313 14231 8347
rect 15577 8313 15611 8347
rect 28457 8313 28491 8347
rect 39957 8313 39991 8347
rect 46857 8313 46891 8347
rect 23765 8245 23799 8279
rect 27445 8245 27479 8279
rect 28273 8245 28307 8279
rect 35265 8245 35299 8279
rect 36277 8245 36311 8279
rect 37289 8245 37323 8279
rect 53481 8245 53515 8279
rect 3249 8041 3283 8075
rect 17509 8041 17543 8075
rect 21557 8041 21591 8075
rect 24593 8041 24627 8075
rect 26065 8041 26099 8075
rect 28641 8041 28675 8075
rect 33057 8041 33091 8075
rect 36461 8041 36495 8075
rect 42257 8041 42291 8075
rect 50169 8041 50203 8075
rect 54033 8041 54067 8075
rect 13001 7973 13035 8007
rect 50537 7973 50571 8007
rect 13369 7905 13403 7939
rect 16221 7905 16255 7939
rect 17693 7905 17727 7939
rect 17785 7905 17819 7939
rect 17969 7905 18003 7939
rect 21557 7905 21591 7939
rect 24501 7905 24535 7939
rect 33609 7905 33643 7939
rect 38761 7905 38795 7939
rect 42809 7905 42843 7939
rect 50629 7905 50663 7939
rect 52653 7905 52687 7939
rect 1869 7837 1903 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4261 7837 4295 7871
rect 6745 7837 6779 7871
rect 7021 7837 7055 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 10793 7837 10827 7871
rect 11621 7837 11655 7871
rect 11805 7837 11839 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 13461 7837 13495 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 16497 7837 16531 7871
rect 17877 7837 17911 7871
rect 19625 7837 19659 7871
rect 21465 7837 21499 7871
rect 24409 7837 24443 7871
rect 26065 7837 26099 7871
rect 26249 7837 26283 7871
rect 26893 7837 26927 7871
rect 27169 7837 27203 7871
rect 27997 7837 28031 7871
rect 28641 7837 28675 7871
rect 28825 7837 28859 7871
rect 36277 7837 36311 7871
rect 38577 7837 38611 7871
rect 50353 7837 50387 7871
rect 2136 7769 2170 7803
rect 3801 7769 3835 7803
rect 19892 7769 19926 7803
rect 27629 7769 27663 7803
rect 27905 7769 27939 7803
rect 33517 7769 33551 7803
rect 42625 7769 42659 7803
rect 52920 7769 52954 7803
rect 6561 7701 6595 7735
rect 6929 7701 6963 7735
rect 11069 7701 11103 7735
rect 11713 7701 11747 7735
rect 21005 7701 21039 7735
rect 21833 7701 21867 7735
rect 24777 7701 24811 7735
rect 26709 7701 26743 7735
rect 27077 7701 27111 7735
rect 27813 7701 27847 7735
rect 28181 7701 28215 7735
rect 33425 7701 33459 7735
rect 42717 7701 42751 7735
rect 1593 7497 1627 7531
rect 2789 7497 2823 7531
rect 13737 7497 13771 7531
rect 17325 7497 17359 7531
rect 20821 7497 20855 7531
rect 35449 7497 35483 7531
rect 36027 7497 36061 7531
rect 53113 7497 53147 7531
rect 16957 7429 16991 7463
rect 17049 7429 17083 7463
rect 24010 7429 24044 7463
rect 27230 7429 27264 7463
rect 32505 7429 32539 7463
rect 35817 7429 35851 7463
rect 37749 7429 37783 7463
rect 43974 7429 44008 7463
rect 1409 7361 1443 7395
rect 2329 7361 2363 7395
rect 2973 7361 3007 7395
rect 6377 7361 6411 7395
rect 6644 7361 6678 7395
rect 9680 7361 9714 7395
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 14105 7361 14139 7395
rect 15301 7361 15335 7395
rect 16681 7361 16715 7395
rect 16829 7361 16863 7395
rect 17146 7361 17180 7395
rect 20545 7361 20579 7395
rect 20637 7361 20671 7395
rect 22477 7361 22511 7395
rect 22753 7361 22787 7395
rect 32321 7361 32355 7395
rect 32413 7361 32447 7395
rect 32643 7361 32677 7395
rect 33609 7361 33643 7395
rect 38577 7361 38611 7395
rect 43729 7361 43763 7395
rect 46397 7361 46431 7395
rect 53021 7361 53055 7395
rect 53205 7361 53239 7395
rect 9413 7293 9447 7327
rect 14197 7293 14231 7327
rect 15577 7293 15611 7327
rect 20821 7293 20855 7327
rect 23765 7293 23799 7327
rect 26985 7293 27019 7327
rect 32781 7293 32815 7327
rect 46673 7293 46707 7327
rect 2145 7225 2179 7259
rect 7757 7225 7791 7259
rect 10793 7225 10827 7259
rect 33793 7225 33827 7259
rect 38761 7225 38795 7259
rect 25145 7157 25179 7191
rect 28365 7157 28399 7191
rect 32137 7157 32171 7191
rect 36001 7157 36035 7191
rect 36185 7157 36219 7191
rect 37841 7157 37875 7191
rect 45109 7157 45143 7191
rect 46213 7157 46247 7191
rect 46581 7157 46615 7191
rect 9781 6953 9815 6987
rect 13553 6953 13587 6987
rect 20361 6953 20395 6987
rect 21557 6953 21591 6987
rect 32873 6953 32907 6987
rect 36001 6953 36035 6987
rect 21005 6885 21039 6919
rect 37197 6885 37231 6919
rect 41889 6885 41923 6919
rect 42349 6885 42383 6919
rect 1685 6817 1719 6851
rect 22201 6817 22235 6851
rect 33517 6817 33551 6851
rect 38301 6817 38335 6851
rect 40877 6817 40911 6851
rect 42809 6817 42843 6851
rect 42901 6817 42935 6851
rect 48953 6817 48987 6851
rect 1409 6749 1443 6783
rect 3157 6749 3191 6783
rect 3801 6749 3835 6783
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 6745 6749 6779 6783
rect 9781 6749 9815 6783
rect 9965 6749 9999 6783
rect 12909 6749 12943 6783
rect 13057 6749 13091 6783
rect 13185 6749 13219 6783
rect 13415 6749 13449 6783
rect 14112 6749 14146 6783
rect 14198 6749 14232 6783
rect 14473 6749 14507 6783
rect 14611 6749 14645 6783
rect 16129 6749 16163 6783
rect 16222 6749 16256 6783
rect 16635 6749 16669 6783
rect 17233 6749 17267 6783
rect 17326 6749 17360 6783
rect 17698 6749 17732 6783
rect 22109 6749 22143 6783
rect 22293 6749 22327 6783
rect 31033 6749 31067 6783
rect 37105 6749 37139 6783
rect 37289 6749 37323 6783
rect 37933 6749 37967 6783
rect 38117 6749 38151 6783
rect 40233 6749 40267 6783
rect 40417 6749 40451 6783
rect 41337 6749 41371 6783
rect 41521 6749 41555 6783
rect 41705 6749 41739 6783
rect 46581 6749 46615 6783
rect 49065 6749 49099 6783
rect 49157 6749 49191 6783
rect 50169 6749 50203 6783
rect 50353 6749 50387 6783
rect 51273 6749 51307 6783
rect 4046 6681 4080 6715
rect 13277 6681 13311 6715
rect 14381 6681 14415 6715
rect 16405 6681 16439 6715
rect 16497 6681 16531 6715
rect 17509 6681 17543 6715
rect 17601 6681 17635 6715
rect 20177 6681 20211 6715
rect 20382 6681 20416 6715
rect 21373 6681 21407 6715
rect 31300 6681 31334 6715
rect 35173 6681 35207 6715
rect 35817 6681 35851 6715
rect 36017 6681 36051 6715
rect 40509 6681 40543 6715
rect 40601 6681 40635 6715
rect 40719 6681 40753 6715
rect 41613 6681 41647 6715
rect 42717 6681 42751 6715
rect 46826 6681 46860 6715
rect 48881 6681 48915 6715
rect 50261 6681 50295 6715
rect 51518 6681 51552 6715
rect 2973 6613 3007 6647
rect 5181 6613 5215 6647
rect 6285 6613 6319 6647
rect 14749 6613 14783 6647
rect 16773 6613 16807 6647
rect 17877 6613 17911 6647
rect 20545 6613 20579 6647
rect 21189 6613 21223 6647
rect 21281 6613 21315 6647
rect 32413 6613 32447 6647
rect 33241 6613 33275 6647
rect 33333 6613 33367 6647
rect 35265 6613 35299 6647
rect 36185 6613 36219 6647
rect 47961 6613 47995 6647
rect 52653 6613 52687 6647
rect 2789 6409 2823 6443
rect 3249 6409 3283 6443
rect 10977 6409 11011 6443
rect 20085 6409 20119 6443
rect 30303 6409 30337 6443
rect 30389 6409 30423 6443
rect 42809 6409 42843 6443
rect 46949 6409 46983 6443
rect 20821 6341 20855 6375
rect 30205 6341 30239 6375
rect 38485 6341 38519 6375
rect 44250 6341 44284 6375
rect 47593 6341 47627 6375
rect 49034 6341 49068 6375
rect 1409 6273 1443 6307
rect 2329 6273 2363 6307
rect 3157 6273 3191 6307
rect 9864 6273 9898 6307
rect 17417 6273 17451 6307
rect 19717 6273 19751 6307
rect 22017 6273 22051 6307
rect 22201 6273 22235 6307
rect 26065 6273 26099 6307
rect 26249 6273 26283 6307
rect 29561 6273 29595 6307
rect 29745 6273 29779 6307
rect 30481 6273 30515 6307
rect 34161 6273 34195 6307
rect 34253 6273 34287 6307
rect 35081 6273 35115 6307
rect 35265 6273 35299 6307
rect 36277 6273 36311 6307
rect 38669 6273 38703 6307
rect 38761 6273 38795 6307
rect 39221 6273 39255 6307
rect 39405 6273 39439 6307
rect 41153 6273 41187 6307
rect 43177 6273 43211 6307
rect 46397 6273 46431 6307
rect 46581 6273 46615 6307
rect 46673 6273 46707 6307
rect 46811 6273 46845 6307
rect 47777 6273 47811 6307
rect 3341 6205 3375 6239
rect 9597 6205 9631 6239
rect 17141 6205 17175 6239
rect 22109 6205 22143 6239
rect 22293 6205 22327 6239
rect 40969 6205 41003 6239
rect 43269 6205 43303 6239
rect 43361 6205 43395 6239
rect 44005 6205 44039 6239
rect 48053 6205 48087 6239
rect 48789 6205 48823 6239
rect 2145 6137 2179 6171
rect 21097 6137 21131 6171
rect 38485 6137 38519 6171
rect 47961 6137 47995 6171
rect 1593 6069 1627 6103
rect 20085 6069 20119 6103
rect 20269 6069 20303 6103
rect 21833 6069 21867 6103
rect 26065 6069 26099 6103
rect 29561 6069 29595 6103
rect 34437 6069 34471 6103
rect 35081 6069 35115 6103
rect 36369 6069 36403 6103
rect 39221 6069 39255 6103
rect 41337 6069 41371 6103
rect 45385 6069 45419 6103
rect 50169 6069 50203 6103
rect 7849 5865 7883 5899
rect 9965 5865 9999 5899
rect 19993 5865 20027 5899
rect 21465 5797 21499 5831
rect 22017 5797 22051 5831
rect 27629 5797 27663 5831
rect 30941 5797 30975 5831
rect 35725 5797 35759 5831
rect 43361 5797 43395 5831
rect 47409 5797 47443 5831
rect 48789 5797 48823 5831
rect 2513 5729 2547 5763
rect 2605 5729 2639 5763
rect 4261 5729 4295 5763
rect 4353 5729 4387 5763
rect 24409 5729 24443 5763
rect 29561 5729 29595 5763
rect 1593 5661 1627 5695
rect 6469 5661 6503 5695
rect 10149 5661 10183 5695
rect 10425 5661 10459 5695
rect 14289 5661 14323 5695
rect 14473 5661 14507 5695
rect 14565 5661 14599 5695
rect 20177 5661 20211 5695
rect 20453 5661 20487 5695
rect 21097 5661 21131 5695
rect 21925 5661 21959 5695
rect 22109 5661 22143 5695
rect 26249 5661 26283 5695
rect 29817 5661 29851 5695
rect 32045 5661 32079 5695
rect 32137 5661 32171 5695
rect 34713 5661 34747 5695
rect 34897 5661 34931 5695
rect 35725 5661 35759 5695
rect 36001 5661 36035 5695
rect 41521 5661 41555 5695
rect 41981 5661 42015 5695
rect 45109 5661 45143 5695
rect 46857 5661 46891 5695
rect 47249 5661 47283 5695
rect 48973 5661 49007 5695
rect 49065 5661 49099 5695
rect 50169 5661 50203 5695
rect 50353 5661 50387 5695
rect 6736 5593 6770 5627
rect 20361 5593 20395 5627
rect 21281 5593 21315 5627
rect 24676 5593 24710 5627
rect 26494 5593 26528 5627
rect 35909 5593 35943 5627
rect 40325 5593 40359 5627
rect 40509 5593 40543 5627
rect 42226 5593 42260 5627
rect 47041 5593 47075 5627
rect 47133 5593 47167 5627
rect 48789 5593 48823 5627
rect 2053 5525 2087 5559
rect 2421 5525 2455 5559
rect 3801 5525 3835 5559
rect 4169 5525 4203 5559
rect 10333 5525 10367 5559
rect 14105 5525 14139 5559
rect 25789 5525 25823 5559
rect 32045 5525 32079 5559
rect 35081 5525 35115 5559
rect 41337 5525 41371 5559
rect 45293 5525 45327 5559
rect 50261 5525 50295 5559
rect 7297 5321 7331 5355
rect 10701 5321 10735 5355
rect 14289 5321 14323 5355
rect 18061 5321 18095 5355
rect 21281 5321 21315 5355
rect 24869 5321 24903 5355
rect 26341 5321 26375 5355
rect 1869 5253 1903 5287
rect 13176 5253 13210 5287
rect 20168 5253 20202 5287
rect 35532 5253 35566 5287
rect 39120 5253 39154 5287
rect 51080 5253 51114 5287
rect 2697 5185 2731 5219
rect 3617 5185 3651 5219
rect 4261 5185 4295 5219
rect 4905 5185 4939 5219
rect 5549 5185 5583 5219
rect 6929 5185 6963 5219
rect 7113 5185 7147 5219
rect 10517 5185 10551 5219
rect 10793 5185 10827 5219
rect 16937 5185 16971 5219
rect 19901 5185 19935 5219
rect 24225 5185 24259 5219
rect 24409 5185 24443 5219
rect 25053 5185 25087 5219
rect 25605 5185 25639 5219
rect 25789 5185 25823 5219
rect 25973 5185 26007 5219
rect 26157 5185 26191 5219
rect 31309 5185 31343 5219
rect 34069 5185 34103 5219
rect 34161 5185 34195 5219
rect 34437 5185 34471 5219
rect 35265 5185 35299 5219
rect 50813 5185 50847 5219
rect 2145 5117 2179 5151
rect 12909 5117 12943 5151
rect 16681 5117 16715 5151
rect 24041 5117 24075 5151
rect 25881 5117 25915 5151
rect 38853 5117 38887 5151
rect 4077 5049 4111 5083
rect 31493 5049 31527 5083
rect 2881 4981 2915 5015
rect 3433 4981 3467 5015
rect 4721 4981 4755 5015
rect 5365 4981 5399 5015
rect 10333 4981 10367 5015
rect 33885 4981 33919 5015
rect 34345 4981 34379 5015
rect 36645 4981 36679 5015
rect 40233 4981 40267 5015
rect 52193 4981 52227 5015
rect 7481 4777 7515 4811
rect 7941 4777 7975 4811
rect 11529 4777 11563 4811
rect 16681 4777 16715 4811
rect 25053 4777 25087 4811
rect 30665 4777 30699 4811
rect 36001 4777 36035 4811
rect 40417 4777 40451 4811
rect 49249 4777 49283 4811
rect 5181 4709 5215 4743
rect 31677 4709 31711 4743
rect 37841 4709 37875 4743
rect 10149 4641 10183 4675
rect 35541 4641 35575 4675
rect 45661 4641 45695 4675
rect 47133 4641 47167 4675
rect 1685 4573 1719 4607
rect 2421 4573 2455 4607
rect 3801 4573 3835 4607
rect 4057 4573 4091 4607
rect 6101 4573 6135 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 10416 4573 10450 4607
rect 15945 4573 15979 4607
rect 16221 4573 16255 4607
rect 16865 4573 16899 4607
rect 17141 4573 17175 4607
rect 19349 4573 19383 4607
rect 24409 4573 24443 4607
rect 24502 4573 24536 4607
rect 24685 4573 24719 4607
rect 24874 4573 24908 4607
rect 27813 4573 27847 4607
rect 30113 4573 30147 4607
rect 30481 4573 30515 4607
rect 31125 4573 31159 4607
rect 31493 4573 31527 4607
rect 33333 4573 33367 4607
rect 33517 4573 33551 4607
rect 33701 4573 33735 4607
rect 35265 4551 35299 4585
rect 35421 4573 35455 4607
rect 35679 4573 35713 4607
rect 35817 4573 35851 4607
rect 37657 4573 37691 4607
rect 39865 4573 39899 4607
rect 40141 4573 40175 4607
rect 40233 4573 40267 4607
rect 46857 4573 46891 4607
rect 48697 4573 48731 4607
rect 48881 4573 48915 4607
rect 49065 4573 49099 4607
rect 6368 4505 6402 4539
rect 16129 4505 16163 4539
rect 17049 4505 17083 4539
rect 19533 4505 19567 4539
rect 24777 4505 24811 4539
rect 27997 4505 28031 4539
rect 30297 4505 30331 4539
rect 30389 4505 30423 4539
rect 31309 4505 31343 4539
rect 31401 4505 31435 4539
rect 33609 4505 33643 4539
rect 40049 4505 40083 4539
rect 40969 4505 41003 4539
rect 45477 4505 45511 4539
rect 48973 4505 49007 4539
rect 1869 4437 1903 4471
rect 2605 4437 2639 4471
rect 15761 4437 15795 4471
rect 19717 4437 19751 4471
rect 33885 4437 33919 4471
rect 41061 4437 41095 4471
rect 3341 4233 3375 4267
rect 3985 4233 4019 4267
rect 5181 4233 5215 4267
rect 6653 4233 6687 4267
rect 6745 4233 6779 4267
rect 7941 4233 7975 4267
rect 14933 4233 14967 4267
rect 31401 4233 31435 4267
rect 43821 4233 43855 4267
rect 13921 4165 13955 4199
rect 45661 4165 45695 4199
rect 46765 4165 46799 4199
rect 47777 4165 47811 4199
rect 48973 4165 49007 4199
rect 2228 4097 2262 4131
rect 3801 4097 3835 4131
rect 5365 4097 5399 4131
rect 6377 4097 6411 4131
rect 6837 4097 6871 4131
rect 7665 4097 7699 4131
rect 8585 4097 8619 4131
rect 9597 4097 9631 4131
rect 10701 4097 10735 4131
rect 12725 4097 12759 4131
rect 15117 4097 15151 4131
rect 16865 4097 16899 4131
rect 19165 4097 19199 4131
rect 22661 4097 22695 4131
rect 23857 4097 23891 4131
rect 25421 4097 25455 4131
rect 25605 4097 25639 4131
rect 25789 4097 25823 4131
rect 25973 4097 26007 4131
rect 28273 4097 28307 4131
rect 28540 4097 28574 4131
rect 30849 4097 30883 4131
rect 31033 4097 31067 4131
rect 31125 4097 31159 4131
rect 31217 4097 31251 4131
rect 32321 4097 32355 4131
rect 37473 4097 37507 4131
rect 38301 4097 38335 4131
rect 38439 4097 38473 4131
rect 38577 4097 38611 4131
rect 38715 4097 38749 4131
rect 40417 4097 40451 4131
rect 41153 4097 41187 4131
rect 41337 4097 41371 4131
rect 41429 4097 41463 4131
rect 41545 4097 41579 4131
rect 42697 4097 42731 4131
rect 45477 4097 45511 4131
rect 45753 4097 45787 4131
rect 45845 4097 45879 4131
rect 46489 4097 46523 4131
rect 46673 4097 46707 4131
rect 46857 4097 46891 4131
rect 47593 4097 47627 4131
rect 47869 4097 47903 4131
rect 47961 4097 47995 4131
rect 48809 4097 48843 4131
rect 49065 4097 49099 4131
rect 49157 4097 49191 4131
rect 1961 4029 1995 4063
rect 7941 4029 7975 4063
rect 12541 4029 12575 4063
rect 22477 4029 22511 4063
rect 25697 4029 25731 4063
rect 37289 4029 37323 4063
rect 42441 4029 42475 4063
rect 8401 3961 8435 3995
rect 10517 3961 10551 3995
rect 23673 3961 23707 3995
rect 41705 3961 41739 3995
rect 46029 3961 46063 3995
rect 48145 3961 48179 3995
rect 49341 3961 49375 3995
rect 4721 3893 4755 3927
rect 7757 3893 7791 3927
rect 9689 3893 9723 3927
rect 12909 3893 12943 3927
rect 16681 3893 16715 3927
rect 18981 3893 19015 3927
rect 22845 3893 22879 3927
rect 26157 3893 26191 3927
rect 29653 3893 29687 3927
rect 32505 3893 32539 3927
rect 37657 3893 37691 3927
rect 38853 3893 38887 3927
rect 40601 3893 40635 3927
rect 47041 3893 47075 3927
rect 2145 3689 2179 3723
rect 5273 3689 5307 3723
rect 7205 3689 7239 3723
rect 9505 3689 9539 3723
rect 36921 3689 36955 3723
rect 38761 3689 38795 3723
rect 42809 3689 42843 3723
rect 47501 3689 47535 3723
rect 12081 3621 12115 3655
rect 16865 3621 16899 3655
rect 23305 3621 23339 3655
rect 4445 3553 4479 3587
rect 13001 3553 13035 3587
rect 15485 3553 15519 3587
rect 25053 3553 25087 3587
rect 36455 3553 36489 3587
rect 57989 3553 58023 3587
rect 1869 3485 1903 3519
rect 2697 3485 2731 3519
rect 3801 3485 3835 3519
rect 4537 3485 4571 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 6653 3485 6687 3519
rect 7389 3485 7423 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 9505 3485 9539 3519
rect 9689 3485 9723 3519
rect 9781 3485 9815 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 12265 3485 12299 3519
rect 12725 3485 12759 3519
rect 14105 3485 14139 3519
rect 14289 3485 14323 3519
rect 15752 3485 15786 3519
rect 17785 3485 17819 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 20453 3485 20487 3519
rect 22661 3485 22695 3519
rect 22754 3485 22788 3519
rect 23029 3485 23063 3519
rect 23167 3485 23201 3519
rect 24685 3485 24719 3519
rect 24873 3485 24907 3519
rect 24970 3485 25004 3519
rect 25248 3485 25282 3519
rect 25881 3485 25915 3519
rect 26148 3485 26182 3519
rect 31033 3485 31067 3519
rect 31309 3485 31343 3519
rect 31401 3485 31435 3519
rect 32137 3485 32171 3519
rect 34897 3485 34931 3519
rect 35173 3485 35207 3519
rect 36185 3485 36219 3519
rect 36357 3485 36391 3519
rect 36599 3485 36633 3519
rect 36737 3485 36771 3519
rect 38209 3485 38243 3519
rect 38577 3485 38611 3519
rect 40509 3485 40543 3519
rect 41245 3485 41279 3519
rect 41521 3485 41555 3519
rect 41613 3485 41647 3519
rect 42257 3485 42291 3519
rect 42529 3485 42563 3519
rect 42625 3485 42659 3519
rect 43269 3485 43303 3519
rect 45201 3485 45235 3519
rect 45937 3485 45971 3519
rect 46121 3485 46155 3519
rect 46305 3485 46339 3519
rect 46949 3485 46983 3519
rect 47133 3485 47167 3519
rect 47363 3485 47397 3519
rect 49065 3485 49099 3519
rect 50169 3485 50203 3519
rect 57713 3485 57747 3519
rect 11437 3417 11471 3451
rect 20720 3417 20754 3451
rect 22937 3417 22971 3451
rect 31217 3417 31251 3451
rect 33517 3417 33551 3451
rect 38393 3417 38427 3451
rect 38485 3417 38519 3451
rect 41429 3417 41463 3451
rect 42441 3417 42475 3451
rect 46213 3417 46247 3451
rect 47225 3417 47259 3451
rect 50414 3417 50448 3451
rect 2881 3349 2915 3383
rect 3985 3349 4019 3383
rect 4629 3349 4663 3383
rect 5825 3349 5859 3383
rect 6469 3349 6503 3383
rect 8217 3349 8251 3383
rect 10977 3349 11011 3383
rect 14473 3349 14507 3383
rect 17969 3349 18003 3383
rect 18521 3349 18555 3383
rect 19257 3349 19291 3383
rect 21833 3349 21867 3383
rect 25421 3349 25455 3383
rect 27261 3349 27295 3383
rect 31585 3349 31619 3383
rect 32229 3349 32263 3383
rect 33609 3349 33643 3383
rect 40693 3349 40727 3383
rect 41797 3349 41831 3383
rect 43453 3349 43487 3383
rect 45385 3349 45419 3383
rect 46489 3349 46523 3383
rect 49249 3349 49283 3383
rect 51549 3349 51583 3383
rect 2145 3145 2179 3179
rect 7297 3145 7331 3179
rect 10517 3145 10551 3179
rect 14105 3145 14139 3179
rect 15853 3145 15887 3179
rect 19717 3145 19751 3179
rect 20453 3145 20487 3179
rect 21097 3145 21131 3179
rect 26985 3145 27019 3179
rect 27629 3145 27663 3179
rect 31493 3145 31527 3179
rect 34805 3145 34839 3179
rect 39589 3145 39623 3179
rect 41337 3145 41371 3179
rect 43821 3145 43855 3179
rect 50537 3145 50571 3179
rect 9404 3077 9438 3111
rect 12909 3077 12943 3111
rect 18604 3077 18638 3111
rect 23029 3077 23063 3111
rect 25136 3077 25170 3111
rect 29368 3077 29402 3111
rect 33692 3077 33726 3111
rect 35532 3077 35566 3111
rect 38476 3077 38510 3111
rect 41061 3077 41095 3111
rect 42686 3077 42720 3111
rect 49402 3077 49436 3111
rect 57161 3077 57195 3111
rect 1869 3009 1903 3043
rect 2697 3009 2731 3043
rect 3433 3009 3467 3043
rect 4712 3009 4746 3043
rect 6377 3009 6411 3043
rect 6561 3009 6595 3043
rect 6745 3009 6779 3043
rect 7481 3009 7515 3043
rect 8677 3009 8711 3043
rect 11713 3009 11747 3043
rect 12541 3009 12575 3043
rect 12725 3009 12759 3043
rect 13921 3009 13955 3043
rect 14749 3009 14783 3043
rect 15393 3009 15427 3043
rect 16037 3009 16071 3043
rect 16865 3009 16899 3043
rect 17601 3009 17635 3043
rect 20637 3009 20671 3043
rect 21281 3009 21315 3043
rect 21833 3009 21867 3043
rect 22661 3009 22695 3043
rect 22754 3009 22788 3043
rect 22937 3009 22971 3043
rect 23167 3009 23201 3043
rect 23765 3009 23799 3043
rect 24869 3009 24903 3043
rect 27169 3009 27203 3043
rect 27813 3009 27847 3043
rect 29101 3009 29135 3043
rect 30941 3009 30975 3043
rect 31125 3009 31159 3043
rect 31217 3009 31251 3043
rect 31309 3009 31343 3043
rect 32413 3009 32447 3043
rect 33425 3009 33459 3043
rect 37289 3009 37323 3043
rect 40049 3009 40083 3043
rect 40785 3009 40819 3043
rect 40969 3009 41003 3043
rect 41153 3009 41187 3043
rect 44281 3009 44315 3043
rect 45661 3009 45695 3043
rect 45928 3009 45962 3043
rect 47593 3009 47627 3043
rect 49157 3009 49191 3043
rect 50997 3009 51031 3043
rect 51733 3009 51767 3043
rect 52929 3009 52963 3043
rect 54401 3009 54435 3043
rect 55873 3009 55907 3043
rect 56885 3009 56919 3043
rect 57897 3009 57931 3043
rect 4445 2941 4479 2975
rect 6837 2941 6871 2975
rect 9137 2941 9171 2975
rect 13737 2941 13771 2975
rect 18337 2941 18371 2975
rect 35265 2941 35299 2975
rect 38209 2941 38243 2975
rect 42441 2941 42475 2975
rect 3617 2873 3651 2907
rect 23949 2873 23983 2907
rect 40233 2873 40267 2907
rect 47777 2873 47811 2907
rect 51181 2873 51215 2907
rect 2881 2805 2915 2839
rect 5825 2805 5859 2839
rect 8493 2805 8527 2839
rect 11529 2805 11563 2839
rect 14565 2805 14599 2839
rect 15209 2805 15243 2839
rect 17049 2805 17083 2839
rect 17785 2805 17819 2839
rect 22017 2805 22051 2839
rect 23305 2805 23339 2839
rect 26249 2805 26283 2839
rect 30481 2805 30515 2839
rect 32597 2805 32631 2839
rect 36645 2805 36679 2839
rect 37473 2805 37507 2839
rect 44465 2805 44499 2839
rect 47041 2805 47075 2839
rect 51917 2805 51951 2839
rect 53113 2805 53147 2839
rect 54585 2805 54619 2839
rect 56057 2805 56091 2839
rect 58081 2805 58115 2839
rect 22753 2601 22787 2635
rect 28825 2601 28859 2635
rect 30297 2601 30331 2635
rect 40417 2601 40451 2635
rect 46029 2601 46063 2635
rect 4721 2533 4755 2567
rect 6561 2533 6595 2567
rect 10609 2533 10643 2567
rect 13185 2533 13219 2567
rect 23397 2533 23431 2567
rect 26065 2533 26099 2567
rect 43085 2533 43119 2567
rect 3249 2465 3283 2499
rect 22385 2465 22419 2499
rect 32413 2465 32447 2499
rect 34713 2465 34747 2499
rect 34989 2465 35023 2499
rect 41245 2465 41279 2499
rect 46765 2465 46799 2499
rect 51273 2465 51307 2499
rect 3801 2397 3835 2431
rect 4537 2397 4571 2431
rect 5549 2397 5583 2431
rect 6377 2397 6411 2431
rect 7113 2397 7147 2431
rect 8953 2397 8987 2431
rect 9689 2397 9723 2431
rect 10425 2397 10459 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13001 2397 13035 2431
rect 14381 2397 14415 2431
rect 15117 2397 15151 2431
rect 15853 2397 15887 2431
rect 17233 2397 17267 2431
rect 17500 2397 17534 2431
rect 19257 2397 19291 2431
rect 19993 2397 20027 2431
rect 20729 2397 20763 2431
rect 22569 2397 22603 2431
rect 23213 2397 23247 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 25881 2397 25915 2431
rect 26985 2397 27019 2431
rect 28089 2397 28123 2431
rect 29009 2397 29043 2431
rect 29561 2397 29595 2431
rect 30481 2397 30515 2431
rect 30941 2397 30975 2431
rect 32137 2397 32171 2431
rect 33885 2397 33919 2431
rect 36001 2397 36035 2431
rect 37289 2397 37323 2431
rect 37565 2397 37599 2431
rect 43913 2397 43947 2431
rect 45477 2397 45511 2431
rect 45661 2397 45695 2431
rect 45845 2397 45879 2431
rect 48789 2397 48823 2431
rect 50169 2397 50203 2431
rect 51089 2397 51123 2431
rect 52745 2397 52779 2431
rect 53941 2397 53975 2431
rect 55321 2397 55355 2431
rect 56793 2397 56827 2431
rect 57897 2397 57931 2431
rect 1501 2329 1535 2363
rect 38669 2329 38703 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 42901 2329 42935 2363
rect 43729 2329 43763 2363
rect 45753 2329 45787 2363
rect 46581 2329 46615 2363
rect 48053 2329 48087 2363
rect 50445 2329 50479 2363
rect 53021 2329 53055 2363
rect 54217 2329 54251 2363
rect 55597 2329 55631 2363
rect 57069 2329 57103 2363
rect 3985 2261 4019 2295
rect 5733 2261 5767 2295
rect 7297 2261 7331 2295
rect 8033 2261 8067 2295
rect 9137 2261 9171 2295
rect 9873 2261 9907 2295
rect 11713 2261 11747 2295
rect 12449 2261 12483 2295
rect 14565 2261 14599 2295
rect 15301 2261 15335 2295
rect 16037 2261 16071 2295
rect 18613 2261 18647 2295
rect 19441 2261 19475 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
rect 24593 2261 24627 2295
rect 25329 2261 25363 2295
rect 27169 2261 27203 2295
rect 28273 2261 28307 2295
rect 29745 2261 29779 2295
rect 31125 2261 31159 2295
rect 34069 2261 34103 2295
rect 36185 2261 36219 2295
rect 38761 2261 38795 2295
rect 48145 2261 48179 2295
rect 48881 2261 48915 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2317 39627 2375 39633
rect 2317 39593 2329 39627
rect 2363 39624 2375 39627
rect 2774 39624 2780 39636
rect 2363 39596 2780 39624
rect 2363 39593 2375 39596
rect 2317 39587 2375 39593
rect 2774 39584 2780 39596
rect 2832 39584 2838 39636
rect 3050 39624 3056 39636
rect 3011 39596 3056 39624
rect 3050 39584 3056 39596
rect 3108 39584 3114 39636
rect 3694 39584 3700 39636
rect 3752 39624 3758 39636
rect 3973 39627 4031 39633
rect 3973 39624 3985 39627
rect 3752 39596 3985 39624
rect 3752 39584 3758 39596
rect 3973 39593 3985 39596
rect 4019 39593 4031 39627
rect 3973 39587 4031 39593
rect 26234 39584 26240 39636
rect 26292 39624 26298 39636
rect 27157 39627 27215 39633
rect 27157 39624 27169 39627
rect 26292 39596 27169 39624
rect 26292 39584 26298 39596
rect 27157 39593 27169 39596
rect 27203 39593 27215 39627
rect 41414 39624 41420 39636
rect 41375 39596 41420 39624
rect 27157 39587 27215 39593
rect 41414 39584 41420 39596
rect 41472 39584 41478 39636
rect 48682 39584 48688 39636
rect 48740 39624 48746 39636
rect 48961 39627 49019 39633
rect 48961 39624 48973 39627
rect 48740 39596 48973 39624
rect 48740 39584 48746 39596
rect 48961 39593 48973 39596
rect 49007 39593 49019 39627
rect 48961 39587 49019 39593
rect 56134 39584 56140 39636
rect 56192 39624 56198 39636
rect 56413 39627 56471 39633
rect 56413 39624 56425 39627
rect 56192 39596 56425 39624
rect 56192 39584 56198 39596
rect 56413 39593 56425 39596
rect 56459 39593 56471 39627
rect 56413 39587 56471 39593
rect 18690 39448 18696 39500
rect 18748 39488 18754 39500
rect 19245 39491 19303 39497
rect 19245 39488 19257 39491
rect 18748 39460 19257 39488
rect 18748 39448 18754 39460
rect 19245 39457 19257 39460
rect 19291 39457 19303 39491
rect 19245 39451 19303 39457
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39420 1455 39423
rect 1762 39420 1768 39432
rect 1443 39392 1768 39420
rect 1443 39389 1455 39392
rect 1397 39383 1455 39389
rect 1762 39380 1768 39392
rect 1820 39380 1826 39432
rect 2133 39423 2191 39429
rect 2133 39389 2145 39423
rect 2179 39420 2191 39423
rect 2314 39420 2320 39432
rect 2179 39392 2320 39420
rect 2179 39389 2191 39392
rect 2133 39383 2191 39389
rect 2314 39380 2320 39392
rect 2372 39380 2378 39432
rect 2866 39420 2872 39432
rect 2827 39392 2872 39420
rect 2866 39380 2872 39392
rect 2924 39380 2930 39432
rect 3789 39423 3847 39429
rect 3789 39389 3801 39423
rect 3835 39420 3847 39423
rect 4062 39420 4068 39432
rect 3835 39392 4068 39420
rect 3835 39389 3847 39392
rect 3789 39383 3847 39389
rect 4062 39380 4068 39392
rect 4120 39380 4126 39432
rect 26973 39423 27031 39429
rect 26973 39389 26985 39423
rect 27019 39420 27031 39423
rect 32122 39420 32128 39432
rect 27019 39392 32128 39420
rect 27019 39389 27031 39392
rect 26973 39383 27031 39389
rect 32122 39380 32128 39392
rect 32180 39380 32186 39432
rect 33686 39380 33692 39432
rect 33744 39420 33750 39432
rect 33781 39423 33839 39429
rect 33781 39420 33793 39423
rect 33744 39392 33793 39420
rect 33744 39380 33750 39392
rect 33781 39389 33793 39392
rect 33827 39389 33839 39423
rect 33781 39383 33839 39389
rect 54754 39380 54760 39432
rect 54812 39420 54818 39432
rect 56229 39423 56287 39429
rect 56229 39420 56241 39423
rect 54812 39392 56241 39420
rect 54812 39380 54818 39392
rect 56229 39389 56241 39392
rect 56275 39389 56287 39423
rect 56229 39383 56287 39389
rect 1578 39284 1584 39296
rect 1539 39256 1584 39284
rect 1578 39244 1584 39256
rect 1636 39244 1642 39296
rect 34057 39287 34115 39293
rect 34057 39253 34069 39287
rect 34103 39284 34115 39287
rect 43438 39284 43444 39296
rect 34103 39256 43444 39284
rect 34103 39253 34115 39256
rect 34057 39247 34115 39253
rect 43438 39244 43444 39256
rect 43496 39244 43502 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 32122 39080 32128 39092
rect 32083 39052 32128 39080
rect 32122 39040 32128 39052
rect 32180 39040 32186 39092
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 13262 38944 13268 38956
rect 1443 38916 13268 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 13262 38904 13268 38916
rect 13320 38904 13326 38956
rect 32309 38947 32367 38953
rect 32309 38913 32321 38947
rect 32355 38944 32367 38947
rect 32490 38944 32496 38956
rect 32355 38916 32496 38944
rect 32355 38913 32367 38916
rect 32309 38907 32367 38913
rect 32490 38904 32496 38916
rect 32548 38904 32554 38956
rect 1578 38740 1584 38752
rect 1539 38712 1584 38740
rect 1578 38700 1584 38712
rect 1636 38700 1642 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1581 38539 1639 38545
rect 1581 38505 1593 38539
rect 1627 38536 1639 38539
rect 2958 38536 2964 38548
rect 1627 38508 2964 38536
rect 1627 38505 1639 38508
rect 1581 38499 1639 38505
rect 2958 38496 2964 38508
rect 3016 38496 3022 38548
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 14458 38332 14464 38344
rect 1443 38304 14464 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 14458 38292 14464 38304
rect 14516 38292 14522 38344
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 1670 37856 1676 37868
rect 1443 37828 1676 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1670 37816 1676 37828
rect 1728 37816 1734 37868
rect 1578 37652 1584 37664
rect 1539 37624 1584 37652
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 12066 36768 12072 36780
rect 1443 36740 12072 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 12066 36728 12072 36740
rect 12124 36728 12130 36780
rect 1578 36632 1584 36644
rect 1539 36604 1584 36632
rect 1578 36592 1584 36604
rect 1636 36592 1642 36644
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 2038 36156 2044 36168
rect 1443 36128 2044 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 2038 36116 2044 36128
rect 2096 36116 2102 36168
rect 1578 36020 1584 36032
rect 1539 35992 1584 36020
rect 1578 35980 1584 35992
rect 1636 35980 1642 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1854 35000 1860 35012
rect 1815 34972 1860 35000
rect 1854 34960 1860 34972
rect 1912 34960 1918 35012
rect 1946 34932 1952 34944
rect 1907 34904 1952 34932
rect 1946 34892 1952 34904
rect 2004 34892 2010 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1578 34728 1584 34740
rect 1539 34700 1584 34728
rect 1578 34688 1584 34700
rect 1636 34688 1642 34740
rect 2133 34731 2191 34737
rect 2133 34697 2145 34731
rect 2179 34728 2191 34731
rect 6546 34728 6552 34740
rect 2179 34700 6552 34728
rect 2179 34697 2191 34700
rect 2133 34691 2191 34697
rect 6546 34688 6552 34700
rect 6604 34688 6610 34740
rect 1397 34595 1455 34601
rect 1397 34561 1409 34595
rect 1443 34561 1455 34595
rect 2314 34592 2320 34604
rect 2275 34564 2320 34592
rect 1397 34555 1455 34561
rect 1412 34524 1440 34555
rect 2314 34552 2320 34564
rect 2372 34552 2378 34604
rect 6178 34524 6184 34536
rect 1412 34496 6184 34524
rect 6178 34484 6184 34496
rect 6236 34484 6242 34536
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 9490 33980 9496 33992
rect 1443 33952 9496 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 9490 33940 9496 33952
rect 9548 33940 9554 33992
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1394 33504 1400 33516
rect 1355 33476 1400 33504
rect 1394 33464 1400 33476
rect 1452 33464 1458 33516
rect 2501 33507 2559 33513
rect 2501 33473 2513 33507
rect 2547 33504 2559 33507
rect 2774 33504 2780 33516
rect 2547 33476 2780 33504
rect 2547 33473 2559 33476
rect 2501 33467 2559 33473
rect 2774 33464 2780 33476
rect 2832 33464 2838 33516
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2222 33436 2228 33448
rect 1719 33408 2228 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2222 33396 2228 33408
rect 2280 33396 2286 33448
rect 2317 33303 2375 33309
rect 2317 33269 2329 33303
rect 2363 33300 2375 33303
rect 6638 33300 6644 33312
rect 2363 33272 6644 33300
rect 2363 33269 2375 33272
rect 2317 33263 2375 33269
rect 6638 33260 6644 33272
rect 6696 33260 6702 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 17034 32892 17040 32904
rect 1443 32864 17040 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32376 1458 32428
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 21910 32212 21916 32224
rect 1627 32184 21916 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 21910 32172 21916 32184
rect 21968 32172 21974 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 2133 32011 2191 32017
rect 2133 31977 2145 32011
rect 2179 32008 2191 32011
rect 4982 32008 4988 32020
rect 2179 31980 4988 32008
rect 2179 31977 2191 31980
rect 2133 31971 2191 31977
rect 4982 31968 4988 31980
rect 5040 31968 5046 32020
rect 15470 31940 15476 31952
rect 1412 31912 15476 31940
rect 1412 31813 1440 31912
rect 15470 31900 15476 31912
rect 15528 31900 15534 31952
rect 1397 31807 1455 31813
rect 1397 31773 1409 31807
rect 1443 31773 1455 31807
rect 2314 31804 2320 31816
rect 2275 31776 2320 31804
rect 1397 31767 1455 31773
rect 2314 31764 2320 31776
rect 2372 31764 2378 31816
rect 1578 31668 1584 31680
rect 1539 31640 1584 31668
rect 1578 31628 1584 31640
rect 1636 31628 1642 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1762 31328 1768 31340
rect 1723 31300 1768 31328
rect 1762 31288 1768 31300
rect 1820 31288 1826 31340
rect 2498 31260 2504 31272
rect 2459 31232 2504 31260
rect 2498 31220 2504 31232
rect 2556 31220 2562 31272
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 12894 30784 12900 30796
rect 1412 30756 12900 30784
rect 1412 30725 1440 30756
rect 12894 30744 12900 30756
rect 12952 30744 12958 30796
rect 1397 30719 1455 30725
rect 1397 30685 1409 30719
rect 1443 30685 1455 30719
rect 2406 30716 2412 30728
rect 2367 30688 2412 30716
rect 1397 30679 1455 30685
rect 2406 30676 2412 30688
rect 2464 30676 2470 30728
rect 3050 30716 3056 30728
rect 3011 30688 3056 30716
rect 3050 30676 3056 30688
rect 3108 30676 3114 30728
rect 4890 30716 4896 30728
rect 4851 30688 4896 30716
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 1578 30580 1584 30592
rect 1539 30552 1584 30580
rect 1578 30540 1584 30552
rect 1636 30540 1642 30592
rect 2225 30583 2283 30589
rect 2225 30549 2237 30583
rect 2271 30580 2283 30583
rect 2314 30580 2320 30592
rect 2271 30552 2320 30580
rect 2271 30549 2283 30552
rect 2225 30543 2283 30549
rect 2314 30540 2320 30552
rect 2372 30540 2378 30592
rect 2682 30540 2688 30592
rect 2740 30580 2746 30592
rect 2869 30583 2927 30589
rect 2869 30580 2881 30583
rect 2740 30552 2881 30580
rect 2740 30540 2746 30552
rect 2869 30549 2881 30552
rect 2915 30549 2927 30583
rect 4706 30580 4712 30592
rect 4667 30552 4712 30580
rect 2869 30543 2927 30549
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 4706 30317 4712 30320
rect 4700 30308 4712 30317
rect 2056 30280 4476 30308
rect 4667 30280 4712 30308
rect 1394 30200 1400 30252
rect 1452 30240 1458 30252
rect 1581 30243 1639 30249
rect 1581 30240 1593 30243
rect 1452 30212 1593 30240
rect 1452 30200 1458 30212
rect 1581 30209 1593 30212
rect 1627 30209 1639 30243
rect 1581 30203 1639 30209
rect 1854 30132 1860 30184
rect 1912 30172 1918 30184
rect 2056 30181 2084 30280
rect 2314 30249 2320 30252
rect 2308 30240 2320 30249
rect 2275 30212 2320 30240
rect 2308 30203 2320 30212
rect 2314 30200 2320 30203
rect 2372 30200 2378 30252
rect 4448 30249 4476 30280
rect 4700 30271 4712 30280
rect 4706 30268 4712 30271
rect 4764 30268 4770 30320
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 2041 30175 2099 30181
rect 2041 30172 2053 30175
rect 1912 30144 2053 30172
rect 1912 30132 1918 30144
rect 2041 30141 2053 30144
rect 2087 30141 2099 30175
rect 2041 30135 2099 30141
rect 1397 30039 1455 30045
rect 1397 30005 1409 30039
rect 1443 30036 1455 30039
rect 3050 30036 3056 30048
rect 1443 30008 3056 30036
rect 1443 30005 1455 30008
rect 1397 29999 1455 30005
rect 3050 29996 3056 30008
rect 3108 29996 3114 30048
rect 3418 30036 3424 30048
rect 3331 30008 3424 30036
rect 3418 29996 3424 30008
rect 3476 30036 3482 30048
rect 5074 30036 5080 30048
rect 3476 30008 5080 30036
rect 3476 29996 3482 30008
rect 5074 29996 5080 30008
rect 5132 29996 5138 30048
rect 5810 30036 5816 30048
rect 5771 30008 5816 30036
rect 5810 29996 5816 30008
rect 5868 29996 5874 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2317 29835 2375 29841
rect 2317 29801 2329 29835
rect 2363 29832 2375 29835
rect 2406 29832 2412 29844
rect 2363 29804 2412 29832
rect 2363 29801 2375 29804
rect 2317 29795 2375 29801
rect 2406 29792 2412 29804
rect 2464 29792 2470 29844
rect 4525 29835 4583 29841
rect 4525 29801 4537 29835
rect 4571 29832 4583 29835
rect 4890 29832 4896 29844
rect 4571 29804 4896 29832
rect 4571 29801 4583 29804
rect 4525 29795 4583 29801
rect 4890 29792 4896 29804
rect 4948 29792 4954 29844
rect 5074 29792 5080 29844
rect 5132 29832 5138 29844
rect 6365 29835 6423 29841
rect 6365 29832 6377 29835
rect 5132 29804 6377 29832
rect 5132 29792 5138 29804
rect 6365 29801 6377 29804
rect 6411 29801 6423 29835
rect 6365 29795 6423 29801
rect 2590 29724 2596 29776
rect 2648 29764 2654 29776
rect 2648 29736 5120 29764
rect 2648 29724 2654 29736
rect 2682 29656 2688 29708
rect 2740 29696 2746 29708
rect 2976 29705 3004 29736
rect 2777 29699 2835 29705
rect 2777 29696 2789 29699
rect 2740 29668 2789 29696
rect 2740 29656 2746 29668
rect 2777 29665 2789 29668
rect 2823 29665 2835 29699
rect 2777 29659 2835 29665
rect 2961 29699 3019 29705
rect 2961 29665 2973 29699
rect 3007 29665 3019 29699
rect 4982 29696 4988 29708
rect 4943 29668 4988 29696
rect 2961 29659 3019 29665
rect 4982 29656 4988 29668
rect 5040 29656 5046 29708
rect 5092 29705 5120 29736
rect 5077 29699 5135 29705
rect 5077 29665 5089 29699
rect 5123 29665 5135 29699
rect 5077 29659 5135 29665
rect 6457 29699 6515 29705
rect 6457 29665 6469 29699
rect 6503 29665 6515 29699
rect 6457 29659 6515 29665
rect 1670 29628 1676 29640
rect 1631 29600 1676 29628
rect 1670 29588 1676 29600
rect 1728 29588 1734 29640
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 5810 29628 5816 29640
rect 4939 29600 5816 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 5810 29588 5816 29600
rect 5868 29628 5874 29640
rect 6472 29628 6500 29659
rect 5868 29600 6500 29628
rect 6641 29631 6699 29637
rect 5868 29588 5874 29600
rect 6641 29597 6653 29631
rect 6687 29628 6699 29631
rect 6730 29628 6736 29640
rect 6687 29600 6736 29628
rect 6687 29597 6699 29600
rect 6641 29591 6699 29597
rect 6730 29588 6736 29600
rect 6788 29588 6794 29640
rect 2685 29563 2743 29569
rect 2685 29529 2697 29563
rect 2731 29560 2743 29563
rect 3418 29560 3424 29572
rect 2731 29532 3424 29560
rect 2731 29529 2743 29532
rect 2685 29523 2743 29529
rect 3418 29520 3424 29532
rect 3476 29520 3482 29572
rect 6362 29560 6368 29572
rect 6323 29532 6368 29560
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 1765 29495 1823 29501
rect 1765 29461 1777 29495
rect 1811 29492 1823 29495
rect 3326 29492 3332 29504
rect 1811 29464 3332 29492
rect 1811 29461 1823 29464
rect 1765 29455 1823 29461
rect 3326 29452 3332 29464
rect 3384 29452 3390 29504
rect 6825 29495 6883 29501
rect 6825 29461 6837 29495
rect 6871 29492 6883 29495
rect 7098 29492 7104 29504
rect 6871 29464 7104 29492
rect 6871 29461 6883 29464
rect 6825 29455 6883 29461
rect 7098 29452 7104 29464
rect 7156 29452 7162 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1670 29248 1676 29300
rect 1728 29288 1734 29300
rect 2130 29288 2136 29300
rect 1728 29260 2136 29288
rect 1728 29248 1734 29260
rect 2130 29248 2136 29260
rect 2188 29248 2194 29300
rect 5629 29291 5687 29297
rect 5629 29257 5641 29291
rect 5675 29257 5687 29291
rect 5629 29251 5687 29257
rect 5644 29220 5672 29251
rect 6362 29248 6368 29300
rect 6420 29288 6426 29300
rect 7745 29291 7803 29297
rect 7745 29288 7757 29291
rect 6420 29260 7757 29288
rect 6420 29248 6426 29260
rect 7745 29257 7757 29260
rect 7791 29257 7803 29291
rect 12894 29288 12900 29300
rect 12855 29260 12900 29288
rect 7745 29251 7803 29257
rect 12894 29248 12900 29260
rect 12952 29248 12958 29300
rect 15470 29288 15476 29300
rect 15431 29260 15476 29288
rect 15470 29248 15476 29260
rect 15528 29248 15534 29300
rect 6610 29223 6668 29229
rect 6610 29220 6622 29223
rect 5644 29192 6622 29220
rect 6610 29189 6622 29192
rect 6656 29189 6668 29223
rect 12342 29220 12348 29232
rect 6610 29183 6668 29189
rect 11532 29192 12348 29220
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29152 1455 29155
rect 2682 29152 2688 29164
rect 1443 29124 2688 29152
rect 1443 29121 1455 29124
rect 1397 29115 1455 29121
rect 2682 29112 2688 29124
rect 2740 29112 2746 29164
rect 2777 29155 2835 29161
rect 2777 29121 2789 29155
rect 2823 29152 2835 29155
rect 2866 29152 2872 29164
rect 2823 29124 2872 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 2866 29112 2872 29124
rect 2924 29112 2930 29164
rect 5810 29152 5816 29164
rect 5771 29124 5816 29152
rect 5810 29112 5816 29124
rect 5868 29112 5874 29164
rect 11532 29161 11560 29192
rect 12342 29180 12348 29192
rect 12400 29220 12406 29232
rect 12400 29192 14136 29220
rect 12400 29180 12406 29192
rect 11517 29155 11575 29161
rect 11517 29121 11529 29155
rect 11563 29121 11575 29155
rect 11517 29115 11575 29121
rect 11784 29155 11842 29161
rect 11784 29121 11796 29155
rect 11830 29152 11842 29155
rect 12158 29152 12164 29164
rect 11830 29124 12164 29152
rect 11830 29121 11842 29124
rect 11784 29115 11842 29121
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 14108 29161 14136 29192
rect 14093 29155 14151 29161
rect 14093 29121 14105 29155
rect 14139 29121 14151 29155
rect 14093 29115 14151 29121
rect 14360 29155 14418 29161
rect 14360 29121 14372 29155
rect 14406 29152 14418 29155
rect 14734 29152 14740 29164
rect 14406 29124 14740 29152
rect 14406 29121 14418 29124
rect 14360 29115 14418 29121
rect 14734 29112 14740 29124
rect 14792 29112 14798 29164
rect 1854 29044 1860 29096
rect 1912 29084 1918 29096
rect 2130 29084 2136 29096
rect 1912 29056 2136 29084
rect 1912 29044 1918 29056
rect 2130 29044 2136 29056
rect 2188 29084 2194 29096
rect 6365 29087 6423 29093
rect 6365 29084 6377 29087
rect 2188 29056 6377 29084
rect 2188 29044 2194 29056
rect 6365 29053 6377 29056
rect 6411 29053 6423 29087
rect 6365 29047 6423 29053
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 2593 29019 2651 29025
rect 2593 28985 2605 29019
rect 2639 29016 2651 29019
rect 2774 29016 2780 29028
rect 2639 28988 2780 29016
rect 2639 28985 2651 28988
rect 2593 28979 2651 28985
rect 2774 28976 2780 28988
rect 2832 28976 2838 29028
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2501 28747 2559 28753
rect 2501 28713 2513 28747
rect 2547 28744 2559 28747
rect 2866 28744 2872 28756
rect 2547 28716 2872 28744
rect 2547 28713 2559 28716
rect 2501 28707 2559 28713
rect 2866 28704 2872 28716
rect 2924 28704 2930 28756
rect 5810 28704 5816 28756
rect 5868 28744 5874 28756
rect 6181 28747 6239 28753
rect 6181 28744 6193 28747
rect 5868 28716 6193 28744
rect 5868 28704 5874 28716
rect 6181 28713 6193 28716
rect 6227 28713 6239 28747
rect 12158 28744 12164 28756
rect 12119 28716 12164 28744
rect 6181 28707 6239 28713
rect 12158 28704 12164 28716
rect 12216 28704 12222 28756
rect 14734 28744 14740 28756
rect 14695 28716 14740 28744
rect 14734 28704 14740 28716
rect 14792 28704 14798 28756
rect 2590 28568 2596 28620
rect 2648 28608 2654 28620
rect 3053 28611 3111 28617
rect 3053 28608 3065 28611
rect 2648 28580 3065 28608
rect 2648 28568 2654 28580
rect 3053 28577 3065 28580
rect 3099 28577 3111 28611
rect 6638 28608 6644 28620
rect 6599 28580 6644 28608
rect 3053 28571 3111 28577
rect 6638 28568 6644 28580
rect 6696 28568 6702 28620
rect 6822 28608 6828 28620
rect 6783 28580 6828 28608
rect 6822 28568 6828 28580
rect 6880 28568 6886 28620
rect 12636 28580 15240 28608
rect 12636 28552 12664 28580
rect 6362 28500 6368 28552
rect 6420 28540 6426 28552
rect 6549 28543 6607 28549
rect 6549 28540 6561 28543
rect 6420 28512 6561 28540
rect 6420 28500 6426 28512
rect 6549 28509 6561 28512
rect 6595 28509 6607 28543
rect 6549 28503 6607 28509
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28509 12403 28543
rect 12618 28540 12624 28552
rect 12579 28512 12624 28540
rect 12345 28503 12403 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 2961 28475 3019 28481
rect 2961 28441 2973 28475
rect 3007 28472 3019 28475
rect 3050 28472 3056 28484
rect 3007 28444 3056 28472
rect 3007 28441 3019 28444
rect 2961 28435 3019 28441
rect 3050 28432 3056 28444
rect 3108 28432 3114 28484
rect 12360 28472 12388 28503
rect 12618 28500 12624 28512
rect 12676 28500 12682 28552
rect 15212 28549 15240 28580
rect 14921 28543 14979 28549
rect 14921 28509 14933 28543
rect 14967 28509 14979 28543
rect 14921 28503 14979 28509
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28540 15255 28543
rect 17126 28540 17132 28552
rect 15243 28512 17132 28540
rect 15243 28509 15255 28512
rect 15197 28503 15255 28509
rect 12529 28475 12587 28481
rect 12360 28444 12434 28472
rect 1762 28364 1768 28416
rect 1820 28404 1826 28416
rect 1949 28407 2007 28413
rect 1949 28404 1961 28407
rect 1820 28376 1961 28404
rect 1820 28364 1826 28376
rect 1949 28373 1961 28376
rect 1995 28373 2007 28407
rect 1949 28367 2007 28373
rect 2869 28407 2927 28413
rect 2869 28373 2881 28407
rect 2915 28404 2927 28407
rect 3878 28404 3884 28416
rect 2915 28376 3884 28404
rect 2915 28373 2927 28376
rect 2869 28367 2927 28373
rect 3878 28364 3884 28376
rect 3936 28364 3942 28416
rect 6730 28364 6736 28416
rect 6788 28404 6794 28416
rect 7282 28404 7288 28416
rect 6788 28376 7288 28404
rect 6788 28364 6794 28376
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 12406 28404 12434 28444
rect 12529 28441 12541 28475
rect 12575 28472 12587 28475
rect 12894 28472 12900 28484
rect 12575 28444 12900 28472
rect 12575 28441 12587 28444
rect 12529 28435 12587 28441
rect 12894 28432 12900 28444
rect 12952 28432 12958 28484
rect 13722 28404 13728 28416
rect 12406 28376 13728 28404
rect 13722 28364 13728 28376
rect 13780 28364 13786 28416
rect 14936 28404 14964 28503
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 17310 28540 17316 28552
rect 17271 28512 17316 28540
rect 17310 28500 17316 28512
rect 17368 28500 17374 28552
rect 15105 28475 15163 28481
rect 15105 28441 15117 28475
rect 15151 28472 15163 28475
rect 15470 28472 15476 28484
rect 15151 28444 15476 28472
rect 15151 28441 15163 28444
rect 15105 28435 15163 28441
rect 15470 28432 15476 28444
rect 15528 28432 15534 28484
rect 17580 28475 17638 28481
rect 17580 28441 17592 28475
rect 17626 28472 17638 28475
rect 18046 28472 18052 28484
rect 17626 28444 18052 28472
rect 17626 28441 17638 28444
rect 17580 28435 17638 28441
rect 18046 28432 18052 28444
rect 18104 28432 18110 28484
rect 16574 28404 16580 28416
rect 14936 28376 16580 28404
rect 16574 28364 16580 28376
rect 16632 28364 16638 28416
rect 18690 28404 18696 28416
rect 18651 28376 18696 28404
rect 18690 28364 18696 28376
rect 18748 28364 18754 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2682 28160 2688 28212
rect 2740 28200 2746 28212
rect 17034 28200 17040 28212
rect 2740 28172 6914 28200
rect 16995 28172 17040 28200
rect 2740 28160 2746 28172
rect 2774 28141 2780 28144
rect 2768 28132 2780 28141
rect 2735 28104 2780 28132
rect 2768 28095 2780 28104
rect 2774 28092 2780 28095
rect 2832 28092 2838 28144
rect 6886 28132 6914 28172
rect 17034 28160 17040 28172
rect 17092 28160 17098 28212
rect 18046 28200 18052 28212
rect 18007 28172 18052 28200
rect 18046 28160 18052 28172
rect 18104 28160 18110 28212
rect 18417 28135 18475 28141
rect 18417 28132 18429 28135
rect 6886 28104 18429 28132
rect 18417 28101 18429 28104
rect 18463 28132 18475 28135
rect 18690 28132 18696 28144
rect 18463 28104 18696 28132
rect 18463 28101 18475 28104
rect 18417 28095 18475 28101
rect 18690 28092 18696 28104
rect 18748 28092 18754 28144
rect 1394 28064 1400 28076
rect 1355 28036 1400 28064
rect 1394 28024 1400 28036
rect 1452 28024 1458 28076
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 17126 28064 17132 28076
rect 17087 28036 17132 28064
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 18230 28064 18236 28076
rect 18191 28036 18236 28064
rect 18230 28024 18236 28036
rect 18288 28024 18294 28076
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 2130 27956 2136 28008
rect 2188 27996 2194 28008
rect 2501 27999 2559 28005
rect 2501 27996 2513 27999
rect 2188 27968 2513 27996
rect 2188 27956 2194 27968
rect 2501 27965 2513 27968
rect 2547 27965 2559 27999
rect 17144 27996 17172 28024
rect 18524 27996 18552 28027
rect 18690 27996 18696 28008
rect 17144 27968 18696 27996
rect 2501 27959 2559 27965
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 3878 27928 3884 27940
rect 3791 27900 3884 27928
rect 3878 27888 3884 27900
rect 3936 27928 3942 27940
rect 6730 27928 6736 27940
rect 3936 27900 6736 27928
rect 3936 27888 3942 27900
rect 6730 27888 6736 27900
rect 6788 27888 6794 27940
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 16666 27860 16672 27872
rect 16627 27832 16672 27860
rect 16666 27820 16672 27832
rect 16724 27820 16730 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 16669 27659 16727 27665
rect 16669 27625 16681 27659
rect 16715 27656 16727 27659
rect 17034 27656 17040 27668
rect 16715 27628 17040 27656
rect 16715 27625 16727 27628
rect 16669 27619 16727 27625
rect 17034 27616 17040 27628
rect 17092 27616 17098 27668
rect 2314 27548 2320 27600
rect 2372 27588 2378 27600
rect 5810 27588 5816 27600
rect 2372 27560 5816 27588
rect 2372 27548 2378 27560
rect 5810 27548 5816 27560
rect 5868 27548 5874 27600
rect 2133 27523 2191 27529
rect 2133 27489 2145 27523
rect 2179 27520 2191 27523
rect 2179 27492 5948 27520
rect 2179 27489 2191 27492
rect 2133 27483 2191 27489
rect 2314 27412 2320 27464
rect 2372 27452 2378 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2372 27424 2881 27452
rect 2372 27412 2378 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 3970 27452 3976 27464
rect 3931 27424 3976 27452
rect 2869 27415 2927 27421
rect 3970 27412 3976 27424
rect 4028 27412 4034 27464
rect 5350 27452 5356 27464
rect 5311 27424 5356 27452
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 5718 27412 5724 27464
rect 5776 27452 5782 27464
rect 5813 27455 5871 27461
rect 5813 27452 5825 27455
rect 5776 27424 5825 27452
rect 5776 27412 5782 27424
rect 5813 27421 5825 27424
rect 5859 27421 5871 27455
rect 5920 27452 5948 27492
rect 6886 27492 10272 27520
rect 6886 27452 6914 27492
rect 5920 27424 6914 27452
rect 5813 27415 5871 27421
rect 9582 27412 9588 27464
rect 9640 27452 9646 27464
rect 10137 27455 10195 27461
rect 10137 27452 10149 27455
rect 9640 27424 10149 27452
rect 9640 27412 9646 27424
rect 10137 27421 10149 27424
rect 10183 27421 10195 27455
rect 10244 27452 10272 27492
rect 12342 27480 12348 27532
rect 12400 27520 12406 27532
rect 15286 27520 15292 27532
rect 12400 27492 15292 27520
rect 12400 27480 12406 27492
rect 15286 27480 15292 27492
rect 15344 27480 15350 27532
rect 15556 27455 15614 27461
rect 10244 27424 11744 27452
rect 10137 27415 10195 27421
rect 1854 27384 1860 27396
rect 1815 27356 1860 27384
rect 1854 27344 1860 27356
rect 1912 27344 1918 27396
rect 6058 27387 6116 27393
rect 6058 27384 6070 27387
rect 5184 27356 6070 27384
rect 2682 27316 2688 27328
rect 2643 27288 2688 27316
rect 2682 27276 2688 27288
rect 2740 27276 2746 27328
rect 2774 27276 2780 27328
rect 2832 27316 2838 27328
rect 5184 27325 5212 27356
rect 6058 27353 6070 27356
rect 6104 27353 6116 27387
rect 6058 27347 6116 27353
rect 6178 27344 6184 27396
rect 6236 27384 6242 27396
rect 10404 27387 10462 27393
rect 6236 27356 10364 27384
rect 6236 27344 6242 27356
rect 3789 27319 3847 27325
rect 3789 27316 3801 27319
rect 2832 27288 3801 27316
rect 2832 27276 2838 27288
rect 3789 27285 3801 27288
rect 3835 27285 3847 27319
rect 3789 27279 3847 27285
rect 5169 27319 5227 27325
rect 5169 27285 5181 27319
rect 5215 27285 5227 27319
rect 5169 27279 5227 27285
rect 6638 27276 6644 27328
rect 6696 27316 6702 27328
rect 7193 27319 7251 27325
rect 7193 27316 7205 27319
rect 6696 27288 7205 27316
rect 6696 27276 6702 27288
rect 7193 27285 7205 27288
rect 7239 27285 7251 27319
rect 10336 27316 10364 27356
rect 10404 27353 10416 27387
rect 10450 27384 10462 27387
rect 10502 27384 10508 27396
rect 10450 27356 10508 27384
rect 10450 27353 10462 27356
rect 10404 27347 10462 27353
rect 10502 27344 10508 27356
rect 10560 27344 10566 27396
rect 10870 27316 10876 27328
rect 10336 27288 10876 27316
rect 7193 27279 7251 27285
rect 10870 27276 10876 27288
rect 10928 27316 10934 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 10928 27288 11529 27316
rect 10928 27276 10934 27288
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 11716 27316 11744 27424
rect 15556 27421 15568 27455
rect 15602 27452 15614 27455
rect 16666 27452 16672 27464
rect 15602 27424 16672 27452
rect 15602 27421 15614 27424
rect 15556 27415 15614 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 25498 27384 25504 27396
rect 12406 27356 25504 27384
rect 12406 27316 12434 27356
rect 25498 27344 25504 27356
rect 25556 27344 25562 27396
rect 11716 27288 12434 27316
rect 11517 27279 11575 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1394 27072 1400 27124
rect 1452 27112 1458 27124
rect 1452 27084 4200 27112
rect 1452 27072 1458 27084
rect 2216 27047 2274 27053
rect 2216 27013 2228 27047
rect 2262 27044 2274 27047
rect 2682 27044 2688 27056
rect 2262 27016 2688 27044
rect 2262 27013 2274 27016
rect 2216 27007 2274 27013
rect 2682 27004 2688 27016
rect 2740 27004 2746 27056
rect 4172 27044 4200 27084
rect 5350 27072 5356 27124
rect 5408 27112 5414 27124
rect 6365 27115 6423 27121
rect 6365 27112 6377 27115
rect 5408 27084 6377 27112
rect 5408 27072 5414 27084
rect 6365 27081 6377 27084
rect 6411 27081 6423 27115
rect 6365 27075 6423 27081
rect 6546 27072 6552 27124
rect 6604 27112 6610 27124
rect 6825 27115 6883 27121
rect 6825 27112 6837 27115
rect 6604 27084 6837 27112
rect 6604 27072 6610 27084
rect 6825 27081 6837 27084
rect 6871 27081 6883 27115
rect 6825 27075 6883 27081
rect 9490 27072 9496 27124
rect 9548 27112 9554 27124
rect 9585 27115 9643 27121
rect 9585 27112 9597 27115
rect 9548 27084 9597 27112
rect 9548 27072 9554 27084
rect 9585 27081 9597 27084
rect 9631 27081 9643 27115
rect 10502 27112 10508 27124
rect 10463 27084 10508 27112
rect 9585 27075 9643 27081
rect 10502 27072 10508 27084
rect 10560 27072 10566 27124
rect 10870 27112 10876 27124
rect 10831 27084 10876 27112
rect 10870 27072 10876 27084
rect 10928 27072 10934 27124
rect 14458 27072 14464 27124
rect 14516 27112 14522 27124
rect 14737 27115 14795 27121
rect 14737 27112 14749 27115
rect 14516 27084 14749 27112
rect 14516 27072 14522 27084
rect 14737 27081 14749 27084
rect 14783 27081 14795 27115
rect 14737 27075 14795 27081
rect 13170 27044 13176 27056
rect 4172 27016 10640 27044
rect 3970 26976 3976 26988
rect 3931 26948 3976 26976
rect 3970 26936 3976 26948
rect 4028 26936 4034 26988
rect 6638 26936 6644 26988
rect 6696 26976 6702 26988
rect 6733 26979 6791 26985
rect 6733 26976 6745 26979
rect 6696 26948 6745 26976
rect 6696 26936 6702 26948
rect 6733 26945 6745 26948
rect 6779 26945 6791 26979
rect 6733 26939 6791 26945
rect 8472 26979 8530 26985
rect 8472 26945 8484 26979
rect 8518 26976 8530 26979
rect 9030 26976 9036 26988
rect 8518 26948 9036 26976
rect 8518 26945 8530 26948
rect 8472 26939 8530 26945
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 1394 26868 1400 26920
rect 1452 26908 1458 26920
rect 1949 26911 2007 26917
rect 1949 26908 1961 26911
rect 1452 26880 1961 26908
rect 1452 26868 1458 26880
rect 1949 26877 1961 26880
rect 1995 26877 2007 26911
rect 1949 26871 2007 26877
rect 1964 26772 1992 26871
rect 6822 26868 6828 26920
rect 6880 26908 6886 26920
rect 6917 26911 6975 26917
rect 6917 26908 6929 26911
rect 6880 26880 6929 26908
rect 6880 26868 6886 26880
rect 6917 26877 6929 26880
rect 6963 26877 6975 26911
rect 6917 26871 6975 26877
rect 8205 26911 8263 26917
rect 8205 26877 8217 26911
rect 8251 26877 8263 26911
rect 8205 26871 8263 26877
rect 3326 26840 3332 26852
rect 3239 26812 3332 26840
rect 3326 26800 3332 26812
rect 3384 26840 3390 26852
rect 5902 26840 5908 26852
rect 3384 26812 5908 26840
rect 3384 26800 3390 26812
rect 5902 26800 5908 26812
rect 5960 26800 5966 26852
rect 2130 26772 2136 26784
rect 1964 26744 2136 26772
rect 2130 26732 2136 26744
rect 2188 26732 2194 26784
rect 3789 26775 3847 26781
rect 3789 26741 3801 26775
rect 3835 26772 3847 26775
rect 4982 26772 4988 26784
rect 3835 26744 4988 26772
rect 3835 26741 3847 26744
rect 3789 26735 3847 26741
rect 4982 26732 4988 26744
rect 5040 26732 5046 26784
rect 6178 26732 6184 26784
rect 6236 26772 6242 26784
rect 8220 26772 8248 26871
rect 6236 26744 8248 26772
rect 10612 26772 10640 27016
rect 10704 27016 13176 27044
rect 10704 26985 10732 27016
rect 13170 27004 13176 27016
rect 13228 27004 13234 27056
rect 10689 26979 10747 26985
rect 10689 26945 10701 26979
rect 10735 26945 10747 26979
rect 10689 26939 10747 26945
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 11020 26948 11065 26976
rect 11020 26936 11026 26948
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 13357 26979 13415 26985
rect 13357 26976 13369 26979
rect 12400 26948 13369 26976
rect 12400 26936 12406 26948
rect 13357 26945 13369 26948
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 13624 26979 13682 26985
rect 13624 26945 13636 26979
rect 13670 26976 13682 26979
rect 14734 26976 14740 26988
rect 13670 26948 14740 26976
rect 13670 26945 13682 26948
rect 13624 26939 13682 26945
rect 14734 26936 14740 26948
rect 14792 26936 14798 26988
rect 15286 26936 15292 26988
rect 15344 26976 15350 26988
rect 17310 26976 17316 26988
rect 15344 26948 17316 26976
rect 15344 26936 15350 26948
rect 17310 26936 17316 26948
rect 17368 26976 17374 26988
rect 18138 26985 18144 26988
rect 17865 26979 17923 26985
rect 17865 26976 17877 26979
rect 17368 26948 17877 26976
rect 17368 26936 17374 26948
rect 17865 26945 17877 26948
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 18132 26939 18144 26985
rect 18196 26976 18202 26988
rect 18196 26948 18232 26976
rect 18138 26936 18144 26939
rect 18196 26936 18202 26948
rect 18598 26772 18604 26784
rect 10612 26744 18604 26772
rect 6236 26732 6242 26744
rect 18598 26732 18604 26744
rect 18656 26772 18662 26784
rect 19245 26775 19303 26781
rect 19245 26772 19257 26775
rect 18656 26744 19257 26772
rect 18656 26732 18662 26744
rect 19245 26741 19257 26744
rect 19291 26741 19303 26775
rect 19245 26735 19303 26741
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2314 26568 2320 26580
rect 2275 26540 2320 26568
rect 2314 26528 2320 26540
rect 2372 26528 2378 26580
rect 5718 26568 5724 26580
rect 5000 26540 5724 26568
rect 2590 26460 2596 26512
rect 2648 26500 2654 26512
rect 4341 26503 4399 26509
rect 2648 26472 2912 26500
rect 2648 26460 2654 26472
rect 2774 26432 2780 26444
rect 2735 26404 2780 26432
rect 2774 26392 2780 26404
rect 2832 26392 2838 26444
rect 2884 26441 2912 26472
rect 4341 26469 4353 26503
rect 4387 26469 4399 26503
rect 4341 26463 4399 26469
rect 2869 26435 2927 26441
rect 2869 26401 2881 26435
rect 2915 26401 2927 26435
rect 4356 26432 4384 26463
rect 5000 26441 5028 26540
rect 5718 26528 5724 26540
rect 5776 26568 5782 26580
rect 6178 26568 6184 26580
rect 5776 26540 6184 26568
rect 5776 26528 5782 26540
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 9030 26528 9036 26580
rect 9088 26568 9094 26580
rect 9125 26571 9183 26577
rect 9125 26568 9137 26571
rect 9088 26540 9137 26568
rect 9088 26528 9094 26540
rect 9125 26537 9137 26540
rect 9171 26537 9183 26571
rect 9125 26531 9183 26537
rect 12437 26571 12495 26577
rect 12437 26537 12449 26571
rect 12483 26568 12495 26571
rect 12618 26568 12624 26580
rect 12483 26540 12624 26568
rect 12483 26537 12495 26540
rect 12437 26531 12495 26537
rect 12618 26528 12624 26540
rect 12676 26528 12682 26580
rect 14734 26568 14740 26580
rect 14695 26540 14740 26568
rect 14734 26528 14740 26540
rect 14792 26528 14798 26580
rect 16758 26568 16764 26580
rect 16132 26540 16764 26568
rect 5994 26460 6000 26512
rect 6052 26500 6058 26512
rect 16132 26500 16160 26540
rect 16758 26528 16764 26540
rect 16816 26568 16822 26580
rect 17497 26571 17555 26577
rect 17497 26568 17509 26571
rect 16816 26540 17509 26568
rect 16816 26528 16822 26540
rect 17497 26537 17509 26540
rect 17543 26537 17555 26571
rect 17497 26531 17555 26537
rect 18138 26528 18144 26580
rect 18196 26568 18202 26580
rect 18233 26571 18291 26577
rect 18233 26568 18245 26571
rect 18196 26540 18245 26568
rect 18196 26528 18202 26540
rect 18233 26537 18245 26540
rect 18279 26537 18291 26571
rect 18233 26531 18291 26537
rect 6052 26472 16160 26500
rect 6052 26460 6058 26472
rect 4985 26435 5043 26441
rect 4356 26404 4844 26432
rect 2869 26395 2927 26401
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26364 1455 26367
rect 4522 26364 4528 26376
rect 1443 26336 4200 26364
rect 4483 26336 4528 26364
rect 1443 26333 1455 26336
rect 1397 26327 1455 26333
rect 2685 26299 2743 26305
rect 2685 26265 2697 26299
rect 2731 26296 2743 26299
rect 3326 26296 3332 26308
rect 2731 26268 3332 26296
rect 2731 26265 2743 26268
rect 2685 26259 2743 26265
rect 3326 26256 3332 26268
rect 3384 26256 3390 26308
rect 4172 26296 4200 26336
rect 4522 26324 4528 26336
rect 4580 26324 4586 26376
rect 4816 26364 4844 26404
rect 4985 26401 4997 26435
rect 5031 26401 5043 26435
rect 13998 26432 14004 26444
rect 4985 26395 5043 26401
rect 6886 26404 14004 26432
rect 5241 26367 5299 26373
rect 5241 26364 5253 26367
rect 4816 26360 4936 26364
rect 5092 26360 5253 26364
rect 4816 26336 5253 26360
rect 4908 26332 5120 26336
rect 5241 26333 5253 26336
rect 5287 26333 5299 26367
rect 5241 26327 5299 26333
rect 6886 26296 6914 26404
rect 13998 26392 14004 26404
rect 14056 26392 14062 26444
rect 14353 26404 14964 26432
rect 9306 26364 9312 26376
rect 9267 26336 9312 26364
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 9490 26364 9496 26376
rect 9451 26336 9496 26364
rect 9490 26324 9496 26336
rect 9548 26324 9554 26376
rect 9585 26367 9643 26373
rect 9585 26333 9597 26367
rect 9631 26364 9643 26367
rect 10134 26364 10140 26376
rect 9631 26336 10140 26364
rect 9631 26333 9643 26336
rect 9585 26327 9643 26333
rect 10134 26324 10140 26336
rect 10192 26364 10198 26376
rect 10962 26364 10968 26376
rect 10192 26336 10968 26364
rect 10192 26324 10198 26336
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 14093 26367 14151 26373
rect 14093 26333 14105 26367
rect 14139 26333 14151 26367
rect 14093 26327 14151 26333
rect 14241 26367 14299 26373
rect 14241 26333 14253 26367
rect 14287 26364 14299 26367
rect 14353 26364 14381 26404
rect 14458 26364 14464 26376
rect 14287 26336 14381 26364
rect 14419 26336 14464 26364
rect 14287 26333 14299 26336
rect 14241 26327 14299 26333
rect 12342 26296 12348 26308
rect 4172 26268 6914 26296
rect 12303 26268 12348 26296
rect 12342 26256 12348 26268
rect 12400 26256 12406 26308
rect 14108 26240 14136 26327
rect 14458 26324 14464 26336
rect 14516 26324 14522 26376
rect 14550 26324 14556 26376
rect 14608 26373 14614 26376
rect 14608 26364 14616 26373
rect 14608 26336 14653 26364
rect 14608 26327 14616 26336
rect 14608 26324 14614 26327
rect 14936 26308 14964 26404
rect 15286 26392 15292 26444
rect 15344 26432 15350 26444
rect 16117 26435 16175 26441
rect 16117 26432 16129 26435
rect 15344 26404 16129 26432
rect 15344 26392 15350 26404
rect 16117 26401 16129 26404
rect 16163 26401 16175 26435
rect 16117 26395 16175 26401
rect 18414 26364 18420 26376
rect 18375 26336 18420 26364
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18598 26364 18604 26376
rect 18559 26336 18604 26364
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 18690 26324 18696 26376
rect 18748 26364 18754 26376
rect 18748 26336 18793 26364
rect 18748 26324 18754 26336
rect 14366 26296 14372 26308
rect 14327 26268 14372 26296
rect 14366 26256 14372 26268
rect 14424 26256 14430 26308
rect 14918 26256 14924 26308
rect 14976 26296 14982 26308
rect 15013 26299 15071 26305
rect 15013 26296 15025 26299
rect 14976 26268 15025 26296
rect 14976 26256 14982 26268
rect 15013 26265 15025 26268
rect 15059 26265 15071 26299
rect 15013 26259 15071 26265
rect 16206 26256 16212 26308
rect 16264 26296 16270 26308
rect 16362 26299 16420 26305
rect 16362 26296 16374 26299
rect 16264 26268 16374 26296
rect 16264 26256 16270 26268
rect 16362 26265 16374 26268
rect 16408 26265 16420 26299
rect 16362 26259 16420 26265
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 6362 26228 6368 26240
rect 6323 26200 6368 26228
rect 6362 26188 6368 26200
rect 6420 26188 6426 26240
rect 14090 26228 14096 26240
rect 14003 26200 14096 26228
rect 14090 26188 14096 26200
rect 14148 26228 14154 26240
rect 15194 26228 15200 26240
rect 14148 26200 15200 26228
rect 14148 26188 14154 26200
rect 15194 26188 15200 26200
rect 15252 26188 15258 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 2590 25984 2596 26036
rect 2648 26024 2654 26036
rect 3973 26027 4031 26033
rect 3973 26024 3985 26027
rect 2648 25996 3985 26024
rect 2648 25984 2654 25996
rect 3973 25993 3985 25996
rect 4019 25993 4031 26027
rect 4522 26024 4528 26036
rect 4483 25996 4528 26024
rect 3973 25987 4031 25993
rect 3988 25956 4016 25987
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 4982 26024 4988 26036
rect 4943 25996 4988 26024
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 16117 26027 16175 26033
rect 16117 25993 16129 26027
rect 16163 26024 16175 26027
rect 16206 26024 16212 26036
rect 16163 25996 16212 26024
rect 16163 25993 16175 25996
rect 16117 25987 16175 25993
rect 16206 25984 16212 25996
rect 16264 25984 16270 26036
rect 4893 25959 4951 25965
rect 3988 25928 4752 25956
rect 1854 25888 1860 25900
rect 1815 25860 1860 25888
rect 1854 25848 1860 25860
rect 1912 25848 1918 25900
rect 2866 25888 2872 25900
rect 2827 25860 2872 25888
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 3881 25891 3939 25897
rect 3881 25857 3893 25891
rect 3927 25888 3939 25891
rect 4614 25888 4620 25900
rect 3927 25860 4620 25888
rect 3927 25857 3939 25860
rect 3881 25851 3939 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 4724 25820 4752 25928
rect 4893 25925 4905 25959
rect 4939 25956 4951 25959
rect 5718 25956 5724 25968
rect 4939 25928 5724 25956
rect 4939 25925 4951 25928
rect 4893 25919 4951 25925
rect 5718 25916 5724 25928
rect 5776 25956 5782 25968
rect 6362 25956 6368 25968
rect 5776 25928 6368 25956
rect 5776 25916 5782 25928
rect 6362 25916 6368 25928
rect 6420 25916 6426 25968
rect 14366 25916 14372 25968
rect 14424 25956 14430 25968
rect 15841 25959 15899 25965
rect 14424 25928 15792 25956
rect 14424 25916 14430 25928
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 12621 25891 12679 25897
rect 12621 25888 12633 25891
rect 12492 25860 12633 25888
rect 12492 25848 12498 25860
rect 12621 25857 12633 25860
rect 12667 25857 12679 25891
rect 12621 25851 12679 25857
rect 12888 25891 12946 25897
rect 12888 25857 12900 25891
rect 12934 25888 12946 25891
rect 14734 25888 14740 25900
rect 12934 25860 14740 25888
rect 12934 25857 12946 25860
rect 12888 25851 12946 25857
rect 14734 25848 14740 25860
rect 14792 25848 14798 25900
rect 15194 25848 15200 25900
rect 15252 25888 15258 25900
rect 15764 25897 15792 25928
rect 15841 25925 15853 25959
rect 15887 25956 15899 25959
rect 16758 25956 16764 25968
rect 15887 25928 16764 25956
rect 15887 25925 15899 25928
rect 15841 25919 15899 25925
rect 16758 25916 16764 25928
rect 16816 25916 16822 25968
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 15252 25860 15485 25888
rect 15252 25848 15258 25860
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 15621 25891 15679 25897
rect 15621 25857 15633 25891
rect 15667 25888 15679 25891
rect 15749 25891 15807 25897
rect 15667 25857 15700 25888
rect 15621 25851 15700 25857
rect 15749 25857 15761 25891
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 5077 25823 5135 25829
rect 5077 25820 5089 25823
rect 4724 25792 5089 25820
rect 5077 25789 5089 25792
rect 5123 25789 5135 25823
rect 15672 25820 15700 25851
rect 15930 25848 15936 25900
rect 15988 25897 15994 25900
rect 15988 25888 15996 25897
rect 15988 25860 16033 25888
rect 15988 25851 15996 25860
rect 15988 25848 15994 25851
rect 16390 25820 16396 25832
rect 15672 25792 16396 25820
rect 5077 25783 5135 25789
rect 16390 25780 16396 25792
rect 16448 25780 16454 25832
rect 2685 25755 2743 25761
rect 2685 25721 2697 25755
rect 2731 25752 2743 25755
rect 5442 25752 5448 25764
rect 2731 25724 5448 25752
rect 2731 25721 2743 25724
rect 2685 25715 2743 25721
rect 5442 25712 5448 25724
rect 5500 25712 5506 25764
rect 2130 25684 2136 25696
rect 2091 25656 2136 25684
rect 2130 25644 2136 25656
rect 2188 25644 2194 25696
rect 2958 25644 2964 25696
rect 3016 25684 3022 25696
rect 14001 25687 14059 25693
rect 14001 25684 14013 25687
rect 3016 25656 14013 25684
rect 3016 25644 3022 25656
rect 14001 25653 14013 25656
rect 14047 25684 14059 25687
rect 14458 25684 14464 25696
rect 14047 25656 14464 25684
rect 14047 25653 14059 25656
rect 14001 25647 14059 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 2130 25440 2136 25492
rect 2188 25480 2194 25492
rect 27062 25480 27068 25492
rect 2188 25452 27068 25480
rect 2188 25440 2194 25452
rect 27062 25440 27068 25452
rect 27120 25440 27126 25492
rect 14734 25412 14740 25424
rect 14695 25384 14740 25412
rect 14734 25372 14740 25384
rect 14792 25372 14798 25424
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25276 1455 25279
rect 2314 25276 2320 25288
rect 1443 25248 2320 25276
rect 1443 25245 1455 25248
rect 1397 25239 1455 25245
rect 2314 25236 2320 25248
rect 2372 25236 2378 25288
rect 2498 25276 2504 25288
rect 2459 25248 2504 25276
rect 2498 25236 2504 25248
rect 2556 25236 2562 25288
rect 5626 25276 5632 25288
rect 5587 25248 5632 25276
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 8846 25236 8852 25288
rect 8904 25276 8910 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8904 25248 8953 25276
rect 8904 25236 8910 25248
rect 8941 25245 8953 25248
rect 8987 25276 8999 25279
rect 9582 25276 9588 25288
rect 8987 25248 9588 25276
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 9582 25236 9588 25248
rect 9640 25276 9646 25288
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 9640 25248 10793 25276
rect 9640 25236 9646 25248
rect 10781 25245 10793 25248
rect 10827 25276 10839 25279
rect 12434 25276 12440 25288
rect 10827 25248 12440 25276
rect 10827 25245 10839 25248
rect 10781 25239 10839 25245
rect 12434 25236 12440 25248
rect 12492 25236 12498 25288
rect 14090 25276 14096 25288
rect 14051 25248 14096 25276
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 14241 25279 14299 25285
rect 14241 25245 14253 25279
rect 14287 25276 14299 25279
rect 14458 25276 14464 25288
rect 14287 25245 14320 25276
rect 14419 25248 14464 25276
rect 14241 25239 14320 25245
rect 4614 25168 4620 25220
rect 4672 25208 4678 25220
rect 6365 25211 6423 25217
rect 6365 25208 6377 25211
rect 4672 25180 6377 25208
rect 4672 25168 4678 25180
rect 6365 25177 6377 25180
rect 6411 25177 6423 25211
rect 6365 25171 6423 25177
rect 9208 25211 9266 25217
rect 9208 25177 9220 25211
rect 9254 25208 9266 25211
rect 10226 25208 10232 25220
rect 9254 25180 10232 25208
rect 9254 25177 9266 25180
rect 9208 25171 9266 25177
rect 10226 25168 10232 25180
rect 10284 25168 10290 25220
rect 11054 25217 11060 25220
rect 11048 25171 11060 25217
rect 11112 25208 11118 25220
rect 11112 25180 11148 25208
rect 11054 25168 11060 25171
rect 11112 25168 11118 25180
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 2317 25143 2375 25149
rect 2317 25109 2329 25143
rect 2363 25140 2375 25143
rect 2406 25140 2412 25152
rect 2363 25112 2412 25140
rect 2363 25109 2375 25112
rect 2317 25103 2375 25109
rect 2406 25100 2412 25112
rect 2464 25100 2470 25152
rect 5445 25143 5503 25149
rect 5445 25109 5457 25143
rect 5491 25140 5503 25143
rect 6270 25140 6276 25152
rect 5491 25112 6276 25140
rect 5491 25109 5503 25112
rect 5445 25103 5503 25109
rect 6270 25100 6276 25112
rect 6328 25100 6334 25152
rect 6641 25143 6699 25149
rect 6641 25109 6653 25143
rect 6687 25140 6699 25143
rect 6822 25140 6828 25152
rect 6687 25112 6828 25140
rect 6687 25109 6699 25112
rect 6641 25103 6699 25109
rect 6822 25100 6828 25112
rect 6880 25140 6886 25152
rect 9858 25140 9864 25152
rect 6880 25112 9864 25140
rect 6880 25100 6886 25112
rect 9858 25100 9864 25112
rect 9916 25100 9922 25152
rect 10042 25100 10048 25152
rect 10100 25140 10106 25152
rect 10321 25143 10379 25149
rect 10321 25140 10333 25143
rect 10100 25112 10333 25140
rect 10100 25100 10106 25112
rect 10321 25109 10333 25112
rect 10367 25109 10379 25143
rect 12158 25140 12164 25152
rect 12119 25112 12164 25140
rect 10321 25103 10379 25109
rect 12158 25100 12164 25112
rect 12216 25100 12222 25152
rect 14292 25140 14320 25239
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 14550 25236 14556 25288
rect 14608 25285 14614 25288
rect 14608 25276 14616 25285
rect 14608 25248 14653 25276
rect 14608 25239 14616 25248
rect 14608 25236 14614 25239
rect 14366 25168 14372 25220
rect 14424 25208 14430 25220
rect 14424 25180 14469 25208
rect 14424 25168 14430 25180
rect 15010 25140 15016 25152
rect 14292 25112 15016 25140
rect 15010 25100 15016 25112
rect 15068 25100 15074 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 5442 24896 5448 24948
rect 5500 24936 5506 24948
rect 5537 24939 5595 24945
rect 5537 24936 5549 24939
rect 5500 24908 5549 24936
rect 5500 24896 5506 24908
rect 5537 24905 5549 24908
rect 5583 24905 5595 24939
rect 5537 24899 5595 24905
rect 10226 24896 10232 24948
rect 10284 24936 10290 24948
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 10284 24908 10333 24936
rect 10284 24896 10290 24908
rect 10321 24905 10333 24908
rect 10367 24905 10379 24939
rect 10321 24899 10379 24905
rect 1670 24828 1676 24880
rect 1728 24868 1734 24880
rect 10042 24868 10048 24880
rect 1728 24840 10048 24868
rect 1728 24828 1734 24840
rect 10042 24828 10048 24840
rect 10100 24828 10106 24880
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 2222 24800 2228 24812
rect 2148 24772 2228 24800
rect 1394 24692 1400 24744
rect 1452 24692 1458 24744
rect 1486 24692 1492 24744
rect 1544 24732 1550 24744
rect 1670 24732 1676 24744
rect 1544 24704 1676 24732
rect 1544 24692 1550 24704
rect 1670 24692 1676 24704
rect 1728 24692 1734 24744
rect 2148 24741 2176 24772
rect 2222 24760 2228 24772
rect 2280 24760 2286 24812
rect 2406 24809 2412 24812
rect 2400 24800 2412 24809
rect 2367 24772 2412 24800
rect 2400 24763 2412 24772
rect 2406 24760 2412 24763
rect 2464 24760 2470 24812
rect 5445 24803 5503 24809
rect 5445 24769 5457 24803
rect 5491 24800 5503 24803
rect 5491 24772 6132 24800
rect 5491 24769 5503 24772
rect 5445 24763 5503 24769
rect 2133 24735 2191 24741
rect 2133 24701 2145 24735
rect 2179 24701 2191 24735
rect 2133 24695 2191 24701
rect 1412 24664 1440 24692
rect 2148 24664 2176 24695
rect 5166 24692 5172 24744
rect 5224 24732 5230 24744
rect 5629 24735 5687 24741
rect 5629 24732 5641 24735
rect 5224 24704 5641 24732
rect 5224 24692 5230 24704
rect 5629 24701 5641 24704
rect 5675 24701 5687 24735
rect 5629 24695 5687 24701
rect 3510 24664 3516 24676
rect 1412 24636 2176 24664
rect 3423 24636 3516 24664
rect 3510 24624 3516 24636
rect 3568 24664 3574 24676
rect 5810 24664 5816 24676
rect 3568 24636 5816 24664
rect 3568 24624 3574 24636
rect 5810 24624 5816 24636
rect 5868 24624 5874 24676
rect 1394 24596 1400 24608
rect 1355 24568 1400 24596
rect 1394 24556 1400 24568
rect 1452 24556 1458 24608
rect 5077 24599 5135 24605
rect 5077 24565 5089 24599
rect 5123 24596 5135 24599
rect 5626 24596 5632 24608
rect 5123 24568 5632 24596
rect 5123 24565 5135 24568
rect 5077 24559 5135 24565
rect 5626 24556 5632 24568
rect 5684 24556 5690 24608
rect 6104 24596 6132 24772
rect 6270 24760 6276 24812
rect 6328 24800 6334 24812
rect 6621 24803 6679 24809
rect 6621 24800 6633 24803
rect 6328 24772 6633 24800
rect 6328 24760 6334 24772
rect 6621 24769 6633 24772
rect 6667 24769 6679 24803
rect 6621 24763 6679 24769
rect 9677 24803 9735 24809
rect 9677 24769 9689 24803
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 6178 24692 6184 24744
rect 6236 24732 6242 24744
rect 6365 24735 6423 24741
rect 6365 24732 6377 24735
rect 6236 24704 6377 24732
rect 6236 24692 6242 24704
rect 6365 24701 6377 24704
rect 6411 24701 6423 24735
rect 9692 24732 9720 24763
rect 9766 24760 9772 24812
rect 9824 24800 9830 24812
rect 9953 24803 10011 24809
rect 9824 24772 9869 24800
rect 9824 24760 9830 24772
rect 9953 24769 9965 24803
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 9968 24732 9996 24763
rect 10134 24760 10140 24812
rect 10192 24809 10198 24812
rect 10192 24800 10200 24809
rect 10192 24772 10237 24800
rect 10192 24763 10200 24772
rect 10192 24760 10198 24763
rect 13630 24760 13636 24812
rect 13688 24800 13694 24812
rect 14550 24800 14556 24812
rect 13688 24772 14556 24800
rect 13688 24760 13694 24772
rect 14550 24760 14556 24772
rect 14608 24800 14614 24812
rect 15654 24800 15660 24812
rect 14608 24772 15660 24800
rect 14608 24760 14614 24772
rect 15654 24760 15660 24772
rect 15712 24800 15718 24812
rect 15930 24800 15936 24812
rect 15712 24772 15936 24800
rect 15712 24760 15718 24772
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 19133 24803 19191 24809
rect 19133 24800 19145 24803
rect 18380 24772 19145 24800
rect 18380 24760 18386 24772
rect 19133 24769 19145 24772
rect 19179 24769 19191 24803
rect 19133 24763 19191 24769
rect 10594 24732 10600 24744
rect 9692 24704 9812 24732
rect 9968 24704 10600 24732
rect 6365 24695 6423 24701
rect 9784 24664 9812 24704
rect 10594 24692 10600 24704
rect 10652 24692 10658 24744
rect 15470 24692 15476 24744
rect 15528 24732 15534 24744
rect 18874 24732 18880 24744
rect 15528 24704 18880 24732
rect 15528 24692 15534 24704
rect 18874 24692 18880 24704
rect 18932 24692 18938 24744
rect 10318 24664 10324 24676
rect 9784 24636 10324 24664
rect 10318 24624 10324 24636
rect 10376 24624 10382 24676
rect 6362 24596 6368 24608
rect 6104 24568 6368 24596
rect 6362 24556 6368 24568
rect 6420 24596 6426 24608
rect 7745 24599 7803 24605
rect 7745 24596 7757 24599
rect 6420 24568 7757 24596
rect 6420 24556 6426 24568
rect 7745 24565 7757 24568
rect 7791 24565 7803 24599
rect 7745 24559 7803 24565
rect 13998 24556 14004 24608
rect 14056 24596 14062 24608
rect 18598 24596 18604 24608
rect 14056 24568 18604 24596
rect 14056 24556 14062 24568
rect 18598 24556 18604 24568
rect 18656 24596 18662 24608
rect 20257 24599 20315 24605
rect 20257 24596 20269 24599
rect 18656 24568 20269 24596
rect 18656 24556 18662 24568
rect 20257 24565 20269 24568
rect 20303 24565 20315 24599
rect 20257 24559 20315 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 2317 24395 2375 24401
rect 2317 24361 2329 24395
rect 2363 24392 2375 24395
rect 2498 24392 2504 24404
rect 2363 24364 2504 24392
rect 2363 24361 2375 24364
rect 2317 24355 2375 24361
rect 2498 24352 2504 24364
rect 2556 24352 2562 24404
rect 6178 24352 6184 24404
rect 6236 24392 6242 24404
rect 8846 24392 8852 24404
rect 6236 24364 8852 24392
rect 6236 24352 6242 24364
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 10965 24395 11023 24401
rect 10965 24361 10977 24395
rect 11011 24392 11023 24395
rect 11054 24392 11060 24404
rect 11011 24364 11060 24392
rect 11011 24361 11023 24364
rect 10965 24355 11023 24361
rect 11054 24352 11060 24364
rect 11112 24352 11118 24404
rect 18233 24395 18291 24401
rect 18233 24361 18245 24395
rect 18279 24392 18291 24395
rect 18322 24392 18328 24404
rect 18279 24364 18328 24392
rect 18279 24361 18291 24364
rect 18233 24355 18291 24361
rect 18322 24352 18328 24364
rect 18380 24352 18386 24404
rect 2406 24284 2412 24336
rect 2464 24324 2470 24336
rect 2464 24296 2912 24324
rect 2464 24284 2470 24296
rect 1394 24216 1400 24268
rect 1452 24256 1458 24268
rect 2884 24265 2912 24296
rect 10318 24284 10324 24336
rect 10376 24324 10382 24336
rect 10376 24296 12434 24324
rect 10376 24284 10382 24296
rect 2777 24259 2835 24265
rect 2777 24256 2789 24259
rect 1452 24228 2789 24256
rect 1452 24216 1458 24228
rect 2777 24225 2789 24228
rect 2823 24225 2835 24259
rect 2777 24219 2835 24225
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 5166 24256 5172 24268
rect 2915 24228 5172 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 5166 24216 5172 24228
rect 5224 24216 5230 24268
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10192 24228 10732 24256
rect 10192 24216 10198 24228
rect 1486 24188 1492 24200
rect 1447 24160 1492 24188
rect 1486 24148 1492 24160
rect 1544 24148 1550 24200
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24188 2743 24191
rect 3510 24188 3516 24200
rect 2731 24160 3516 24188
rect 2731 24157 2743 24160
rect 2685 24151 2743 24157
rect 3510 24148 3516 24160
rect 3568 24148 3574 24200
rect 10226 24188 10232 24200
rect 3620 24160 10232 24188
rect 1670 24080 1676 24132
rect 1728 24120 1734 24132
rect 3620 24120 3648 24160
rect 10226 24148 10232 24160
rect 10284 24148 10290 24200
rect 10318 24148 10324 24200
rect 10376 24188 10382 24200
rect 10502 24197 10508 24200
rect 10469 24191 10508 24197
rect 10376 24160 10421 24188
rect 10376 24148 10382 24160
rect 10469 24157 10481 24191
rect 10469 24151 10508 24157
rect 10502 24148 10508 24151
rect 10560 24148 10566 24200
rect 10704 24188 10732 24228
rect 10786 24191 10844 24197
rect 10786 24188 10798 24191
rect 10704 24160 10798 24188
rect 10786 24157 10798 24160
rect 10832 24157 10844 24191
rect 12406 24188 12434 24296
rect 12526 24216 12532 24268
rect 12584 24256 12590 24268
rect 15470 24256 15476 24268
rect 12584 24228 15476 24256
rect 12584 24216 12590 24228
rect 15470 24216 15476 24228
rect 15528 24256 15534 24268
rect 15565 24259 15623 24265
rect 15565 24256 15577 24259
rect 15528 24228 15577 24256
rect 15528 24216 15534 24228
rect 15565 24225 15577 24228
rect 15611 24225 15623 24259
rect 15565 24219 15623 24225
rect 18874 24216 18880 24268
rect 18932 24256 18938 24268
rect 19245 24259 19303 24265
rect 19245 24256 19257 24259
rect 18932 24228 19257 24256
rect 18932 24216 18938 24228
rect 19245 24225 19257 24228
rect 19291 24225 19303 24259
rect 19245 24219 19303 24225
rect 12710 24188 12716 24200
rect 12406 24160 12716 24188
rect 10786 24151 10844 24157
rect 12710 24148 12716 24160
rect 12768 24188 12774 24200
rect 12897 24191 12955 24197
rect 12897 24188 12909 24191
rect 12768 24160 12909 24188
rect 12768 24148 12774 24160
rect 12897 24157 12909 24160
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 12990 24191 13048 24197
rect 12990 24157 13002 24191
rect 13036 24157 13048 24191
rect 13262 24188 13268 24200
rect 13223 24160 13268 24188
rect 12990 24151 13048 24157
rect 1728 24092 3648 24120
rect 1728 24080 1734 24092
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 4985 24123 5043 24129
rect 4985 24120 4997 24123
rect 4672 24092 4997 24120
rect 4672 24080 4678 24092
rect 4985 24089 4997 24092
rect 5031 24089 5043 24123
rect 10594 24120 10600 24132
rect 10555 24092 10600 24120
rect 4985 24083 5043 24089
rect 10594 24080 10600 24092
rect 10652 24080 10658 24132
rect 10689 24123 10747 24129
rect 10689 24089 10701 24123
rect 10735 24120 10747 24123
rect 12158 24120 12164 24132
rect 10735 24092 12164 24120
rect 10735 24089 10747 24092
rect 10689 24083 10747 24089
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 12802 24080 12808 24132
rect 12860 24120 12866 24132
rect 13004 24120 13032 24151
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 13403 24191 13461 24197
rect 13403 24157 13415 24191
rect 13449 24188 13461 24191
rect 13630 24188 13636 24200
rect 13449 24160 13636 24188
rect 13449 24157 13461 24160
rect 13403 24151 13461 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24188 18475 24191
rect 18690 24188 18696 24200
rect 18463 24160 18552 24188
rect 18651 24160 18696 24188
rect 18463 24157 18475 24160
rect 18417 24151 18475 24157
rect 12860 24092 13032 24120
rect 13173 24123 13231 24129
rect 12860 24080 12866 24092
rect 13173 24089 13185 24123
rect 13219 24120 13231 24123
rect 14366 24120 14372 24132
rect 13219 24092 14372 24120
rect 13219 24089 13231 24092
rect 13173 24083 13231 24089
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 15838 24129 15844 24132
rect 15832 24083 15844 24129
rect 15896 24120 15902 24132
rect 15896 24092 15932 24120
rect 15838 24080 15844 24083
rect 15896 24080 15902 24092
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 2038 24012 2044 24064
rect 2096 24052 2102 24064
rect 13354 24052 13360 24064
rect 2096 24024 13360 24052
rect 2096 24012 2102 24024
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 13538 24052 13544 24064
rect 13499 24024 13544 24052
rect 13538 24012 13544 24024
rect 13596 24012 13602 24064
rect 16942 24052 16948 24064
rect 16903 24024 16948 24052
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 18524 24052 18552 24160
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 18598 24080 18604 24132
rect 18656 24120 18662 24132
rect 18656 24092 18701 24120
rect 18656 24080 18662 24092
rect 19058 24080 19064 24132
rect 19116 24120 19122 24132
rect 19490 24123 19548 24129
rect 19490 24120 19502 24123
rect 19116 24092 19502 24120
rect 19116 24080 19122 24092
rect 19490 24089 19502 24092
rect 19536 24089 19548 24123
rect 19490 24083 19548 24089
rect 20254 24052 20260 24064
rect 18524 24024 20260 24052
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 20622 24052 20628 24064
rect 20583 24024 20628 24052
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 2314 23808 2320 23860
rect 2372 23848 2378 23860
rect 2372 23820 12434 23848
rect 2372 23808 2378 23820
rect 2590 23780 2596 23792
rect 1412 23752 2596 23780
rect 1412 23721 1440 23752
rect 2590 23740 2596 23752
rect 2648 23740 2654 23792
rect 6362 23780 6368 23792
rect 6323 23752 6368 23780
rect 6362 23740 6368 23752
rect 6420 23780 6426 23792
rect 6914 23780 6920 23792
rect 6420 23752 6920 23780
rect 6420 23740 6426 23752
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 12161 23783 12219 23789
rect 12161 23780 12173 23783
rect 10192 23752 12173 23780
rect 10192 23740 10198 23752
rect 12161 23749 12173 23752
rect 12207 23749 12219 23783
rect 12161 23743 12219 23749
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23712 2191 23715
rect 2222 23712 2228 23724
rect 2179 23684 2228 23712
rect 2179 23681 2191 23684
rect 2133 23675 2191 23681
rect 2222 23672 2228 23684
rect 2280 23672 2286 23724
rect 2400 23715 2458 23721
rect 2400 23681 2412 23715
rect 2446 23712 2458 23715
rect 2682 23712 2688 23724
rect 2446 23684 2688 23712
rect 2446 23681 2458 23684
rect 2400 23675 2458 23681
rect 2682 23672 2688 23684
rect 2740 23672 2746 23724
rect 5074 23672 5080 23724
rect 5132 23712 5138 23724
rect 6641 23715 6699 23721
rect 6641 23712 6653 23715
rect 5132 23684 6653 23712
rect 5132 23672 5138 23684
rect 6641 23681 6653 23684
rect 6687 23712 6699 23715
rect 7190 23712 7196 23724
rect 6687 23684 7196 23712
rect 6687 23681 6699 23684
rect 6641 23675 6699 23681
rect 7190 23672 7196 23684
rect 7248 23672 7254 23724
rect 9116 23715 9174 23721
rect 9116 23681 9128 23715
rect 9162 23712 9174 23715
rect 10410 23712 10416 23724
rect 9162 23684 10416 23712
rect 9162 23681 9174 23684
rect 9116 23675 9174 23681
rect 10410 23672 10416 23684
rect 10468 23672 10474 23724
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23712 12035 23715
rect 12066 23712 12072 23724
rect 12023 23684 12072 23712
rect 12023 23681 12035 23684
rect 11977 23675 12035 23681
rect 12066 23672 12072 23684
rect 12124 23672 12130 23724
rect 12406 23712 12434 23820
rect 13354 23808 13360 23860
rect 13412 23848 13418 23860
rect 15838 23848 15844 23860
rect 13412 23820 15700 23848
rect 15799 23820 15844 23848
rect 13412 23808 13418 23820
rect 13072 23783 13130 23789
rect 13072 23749 13084 23783
rect 13118 23780 13130 23783
rect 13538 23780 13544 23792
rect 13118 23752 13544 23780
rect 13118 23749 13130 23752
rect 13072 23743 13130 23749
rect 13538 23740 13544 23752
rect 13596 23740 13602 23792
rect 14366 23740 14372 23792
rect 14424 23780 14430 23792
rect 14826 23780 14832 23792
rect 14424 23752 14832 23780
rect 14424 23740 14430 23752
rect 14826 23740 14832 23752
rect 14884 23780 14890 23792
rect 15473 23783 15531 23789
rect 15473 23780 15485 23783
rect 14884 23752 15485 23780
rect 14884 23740 14890 23752
rect 15473 23749 15485 23752
rect 15519 23749 15531 23783
rect 15473 23743 15531 23749
rect 15565 23783 15623 23789
rect 15565 23749 15577 23783
rect 15611 23780 15623 23783
rect 15672 23780 15700 23820
rect 15838 23808 15844 23820
rect 15896 23808 15902 23860
rect 19058 23848 19064 23860
rect 19019 23820 19064 23848
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 20530 23848 20536 23860
rect 19260 23820 20536 23848
rect 16942 23780 16948 23792
rect 15611 23752 16948 23780
rect 15611 23749 15623 23752
rect 15565 23743 15623 23749
rect 16942 23740 16948 23752
rect 17000 23740 17006 23792
rect 12406 23684 15148 23712
rect 5810 23604 5816 23656
rect 5868 23644 5874 23656
rect 6457 23647 6515 23653
rect 6457 23644 6469 23647
rect 5868 23616 6469 23644
rect 5868 23604 5874 23616
rect 6457 23613 6469 23616
rect 6503 23613 6515 23647
rect 8846 23644 8852 23656
rect 8759 23616 8852 23644
rect 6457 23607 6515 23613
rect 8846 23604 8852 23616
rect 8904 23604 8910 23656
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12492 23616 12817 23644
rect 12492 23604 12498 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 12805 23607 12863 23613
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 2038 23508 2044 23520
rect 1820 23480 2044 23508
rect 1820 23468 1826 23480
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 3510 23508 3516 23520
rect 3471 23480 3516 23508
rect 3510 23468 3516 23480
rect 3568 23468 3574 23520
rect 6362 23508 6368 23520
rect 6323 23480 6368 23508
rect 6362 23468 6368 23480
rect 6420 23468 6426 23520
rect 6825 23511 6883 23517
rect 6825 23477 6837 23511
rect 6871 23508 6883 23511
rect 7466 23508 7472 23520
rect 6871 23480 7472 23508
rect 6871 23477 6883 23480
rect 6825 23471 6883 23477
rect 7466 23468 7472 23480
rect 7524 23468 7530 23520
rect 8864 23508 8892 23604
rect 10226 23576 10232 23588
rect 10187 23548 10232 23576
rect 10226 23536 10232 23548
rect 10284 23536 10290 23588
rect 9582 23508 9588 23520
rect 8864 23480 9588 23508
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 12820 23508 12848 23607
rect 15120 23576 15148 23684
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15345 23715 15403 23721
rect 15252 23684 15297 23712
rect 15252 23672 15258 23684
rect 15345 23681 15357 23715
rect 15391 23712 15403 23715
rect 15391 23681 15424 23712
rect 15345 23675 15424 23681
rect 15396 23644 15424 23675
rect 15654 23672 15660 23724
rect 15712 23721 15718 23724
rect 19260 23721 19288 23820
rect 20530 23808 20536 23820
rect 20588 23808 20594 23860
rect 20622 23780 20628 23792
rect 19444 23752 20628 23780
rect 19444 23721 19472 23752
rect 20622 23740 20628 23752
rect 20680 23740 20686 23792
rect 15712 23712 15720 23721
rect 19245 23715 19303 23721
rect 15712 23684 15757 23712
rect 15712 23675 15720 23684
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23681 19579 23715
rect 19521 23675 19579 23681
rect 15712 23672 15718 23675
rect 16482 23644 16488 23656
rect 15396 23616 16488 23644
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 19444 23576 19472 23675
rect 15120 23548 19472 23576
rect 12986 23508 12992 23520
rect 12820 23480 12992 23508
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13446 23468 13452 23520
rect 13504 23508 13510 23520
rect 14185 23511 14243 23517
rect 14185 23508 14197 23511
rect 13504 23480 14197 23508
rect 13504 23468 13510 23480
rect 14185 23477 14197 23480
rect 14231 23477 14243 23511
rect 14185 23471 14243 23477
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15746 23508 15752 23520
rect 15252 23480 15752 23508
rect 15252 23468 15258 23480
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 19536 23508 19564 23675
rect 18748 23480 19564 23508
rect 18748 23468 18754 23480
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 2682 23304 2688 23316
rect 2643 23276 2688 23304
rect 2682 23264 2688 23276
rect 2740 23264 2746 23316
rect 5810 23304 5816 23316
rect 5771 23276 5816 23304
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 6457 23307 6515 23313
rect 6457 23304 6469 23307
rect 5960 23276 6469 23304
rect 5960 23264 5966 23276
rect 6457 23273 6469 23276
rect 6503 23273 6515 23307
rect 10410 23304 10416 23316
rect 10371 23276 10416 23304
rect 6457 23267 6515 23273
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 14826 23304 14832 23316
rect 14787 23276 14832 23304
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 5997 23239 6055 23245
rect 5997 23205 6009 23239
rect 6043 23236 6055 23239
rect 7650 23236 7656 23248
rect 6043 23208 7656 23236
rect 6043 23205 6055 23208
rect 5997 23199 6055 23205
rect 7650 23196 7656 23208
rect 7708 23196 7714 23248
rect 10318 23236 10324 23248
rect 9784 23208 10324 23236
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 5718 23168 5724 23180
rect 5679 23140 5724 23168
rect 5718 23128 5724 23140
rect 5776 23168 5782 23180
rect 6638 23168 6644 23180
rect 5776 23140 6500 23168
rect 6599 23140 6644 23168
rect 5776 23128 5782 23140
rect 1670 23100 1676 23112
rect 1631 23072 1676 23100
rect 1670 23060 1676 23072
rect 1728 23060 1734 23112
rect 2222 23060 2228 23112
rect 2280 23100 2286 23112
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2280 23072 2881 23100
rect 2280 23060 2286 23072
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 3970 23100 3976 23112
rect 3931 23072 3976 23100
rect 2869 23063 2927 23069
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 5813 23103 5871 23109
rect 5813 23100 5825 23103
rect 4632 23072 5825 23100
rect 3510 22992 3516 23044
rect 3568 23032 3574 23044
rect 4632 23032 4660 23072
rect 5813 23069 5825 23072
rect 5859 23100 5871 23103
rect 6362 23100 6368 23112
rect 5859 23072 6368 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6362 23060 6368 23072
rect 6420 23060 6426 23112
rect 6472 23100 6500 23140
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 9784 23109 9812 23208
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 13449 23239 13507 23245
rect 13449 23205 13461 23239
rect 13495 23236 13507 23239
rect 13630 23236 13636 23248
rect 13495 23208 13636 23236
rect 13495 23205 13507 23208
rect 13449 23199 13507 23205
rect 13630 23196 13636 23208
rect 13688 23196 13694 23248
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 10100 23140 10272 23168
rect 10100 23128 10106 23140
rect 9950 23109 9956 23112
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6472 23072 6745 23100
rect 6733 23069 6745 23072
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 9769 23103 9827 23109
rect 9769 23069 9781 23103
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 9917 23103 9956 23109
rect 9917 23069 9929 23103
rect 9917 23063 9956 23069
rect 9950 23060 9956 23063
rect 10008 23060 10014 23112
rect 10134 23100 10140 23112
rect 10095 23072 10140 23100
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 10244 23109 10272 23140
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 16025 23171 16083 23177
rect 16025 23168 16037 23171
rect 15528 23140 16037 23168
rect 15528 23128 15534 23140
rect 16025 23137 16037 23140
rect 16071 23137 16083 23171
rect 16025 23131 16083 23137
rect 10234 23103 10292 23109
rect 10234 23069 10246 23103
rect 10280 23069 10292 23103
rect 10234 23063 10292 23069
rect 11701 23103 11759 23109
rect 11701 23069 11713 23103
rect 11747 23100 11759 23103
rect 12066 23100 12072 23112
rect 11747 23072 12072 23100
rect 11747 23069 11759 23072
rect 11701 23063 11759 23069
rect 12066 23060 12072 23072
rect 12124 23100 12130 23112
rect 13265 23103 13323 23109
rect 13265 23100 13277 23103
rect 12124 23072 13277 23100
rect 12124 23060 12130 23072
rect 13265 23069 13277 23072
rect 13311 23069 13323 23103
rect 13265 23063 13323 23069
rect 14737 23103 14795 23109
rect 14737 23069 14749 23103
rect 14783 23100 14795 23103
rect 14826 23100 14832 23112
rect 14783 23072 14832 23100
rect 14783 23069 14795 23072
rect 14737 23063 14795 23069
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 21729 23103 21787 23109
rect 21729 23100 21741 23103
rect 21692 23072 21741 23100
rect 21692 23060 21698 23072
rect 21729 23069 21741 23072
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 24670 23060 24676 23112
rect 24728 23100 24734 23112
rect 25409 23103 25467 23109
rect 25409 23100 25421 23103
rect 24728 23072 25421 23100
rect 24728 23060 24734 23072
rect 25409 23069 25421 23072
rect 25455 23069 25467 23103
rect 25409 23063 25467 23069
rect 27982 23060 27988 23112
rect 28040 23100 28046 23112
rect 28629 23103 28687 23109
rect 28629 23100 28641 23103
rect 28040 23072 28641 23100
rect 28040 23060 28046 23072
rect 28629 23069 28641 23072
rect 28675 23069 28687 23103
rect 31202 23100 31208 23112
rect 31163 23072 31208 23100
rect 28629 23063 28687 23069
rect 31202 23060 31208 23072
rect 31260 23100 31266 23112
rect 34606 23100 34612 23112
rect 31260 23072 34612 23100
rect 31260 23060 31266 23072
rect 34606 23060 34612 23072
rect 34664 23060 34670 23112
rect 3568 23004 4660 23032
rect 5537 23035 5595 23041
rect 3568 22992 3574 23004
rect 5537 23001 5549 23035
rect 5583 23032 5595 23035
rect 5902 23032 5908 23044
rect 5583 23004 5908 23032
rect 5583 23001 5595 23004
rect 5537 22995 5595 23001
rect 5902 22992 5908 23004
rect 5960 22992 5966 23044
rect 6457 23035 6515 23041
rect 6457 23001 6469 23035
rect 6503 23032 6515 23035
rect 7834 23032 7840 23044
rect 6503 23004 7840 23032
rect 6503 23001 6515 23004
rect 6457 22995 6515 23001
rect 7834 22992 7840 23004
rect 7892 22992 7898 23044
rect 10045 23035 10103 23041
rect 10045 23001 10057 23035
rect 10091 23032 10103 23035
rect 10318 23032 10324 23044
rect 10091 23004 10324 23032
rect 10091 23001 10103 23004
rect 10045 22995 10103 23001
rect 10318 22992 10324 23004
rect 10376 23032 10382 23044
rect 10594 23032 10600 23044
rect 10376 23004 10600 23032
rect 10376 22992 10382 23004
rect 10594 22992 10600 23004
rect 10652 22992 10658 23044
rect 12529 23035 12587 23041
rect 12529 23032 12541 23035
rect 12406 23004 12541 23032
rect 12406 22976 12434 23004
rect 12529 23001 12541 23004
rect 12575 23001 12587 23035
rect 12529 22995 12587 23001
rect 12713 23035 12771 23041
rect 12713 23001 12725 23035
rect 12759 23032 12771 23035
rect 12894 23032 12900 23044
rect 12759 23004 12900 23032
rect 12759 23001 12771 23004
rect 12713 22995 12771 23001
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 16292 23035 16350 23041
rect 16292 23001 16304 23035
rect 16338 23032 16350 23035
rect 16758 23032 16764 23044
rect 16338 23004 16764 23032
rect 16338 23001 16350 23004
rect 16292 22995 16350 23001
rect 16758 22992 16764 23004
rect 16816 22992 16822 23044
rect 21996 23035 22054 23041
rect 21996 23001 22008 23035
rect 22042 23032 22054 23035
rect 22094 23032 22100 23044
rect 22042 23004 22100 23032
rect 22042 23001 22054 23004
rect 21996 22995 22054 23001
rect 22094 22992 22100 23004
rect 22152 22992 22158 23044
rect 25676 23035 25734 23041
rect 25676 23001 25688 23035
rect 25722 23032 25734 23035
rect 25774 23032 25780 23044
rect 25722 23004 25780 23032
rect 25722 23001 25734 23004
rect 25676 22995 25734 23001
rect 25774 22992 25780 23004
rect 25832 22992 25838 23044
rect 31478 23041 31484 23044
rect 31472 22995 31484 23041
rect 31536 23032 31542 23044
rect 31536 23004 31572 23032
rect 31478 22992 31484 22995
rect 31536 22992 31542 23004
rect 2682 22924 2688 22976
rect 2740 22964 2746 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 2740 22936 3801 22964
rect 2740 22924 2746 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7374 22964 7380 22976
rect 6963 22936 7380 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7374 22924 7380 22936
rect 7432 22924 7438 22976
rect 11882 22964 11888 22976
rect 11843 22936 11888 22964
rect 11882 22924 11888 22936
rect 11940 22964 11946 22976
rect 12342 22964 12348 22976
rect 11940 22936 12348 22964
rect 11940 22924 11946 22936
rect 12342 22924 12348 22936
rect 12400 22936 12434 22976
rect 17402 22964 17408 22976
rect 17363 22936 17408 22964
rect 12400 22924 12406 22936
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 21726 22924 21732 22976
rect 21784 22964 21790 22976
rect 23109 22967 23167 22973
rect 23109 22964 23121 22967
rect 21784 22936 23121 22964
rect 21784 22924 21790 22936
rect 23109 22933 23121 22936
rect 23155 22933 23167 22967
rect 26786 22964 26792 22976
rect 26747 22936 26792 22964
rect 23109 22927 23167 22933
rect 26786 22924 26792 22936
rect 26844 22924 26850 22976
rect 28442 22964 28448 22976
rect 28403 22936 28448 22964
rect 28442 22924 28448 22936
rect 28500 22924 28506 22976
rect 32214 22924 32220 22976
rect 32272 22964 32278 22976
rect 32585 22967 32643 22973
rect 32585 22964 32597 22967
rect 32272 22936 32597 22964
rect 32272 22924 32278 22936
rect 32585 22933 32597 22936
rect 32631 22933 32643 22967
rect 32585 22927 32643 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 2222 22760 2228 22772
rect 2183 22732 2228 22760
rect 2222 22720 2228 22732
rect 2280 22720 2286 22772
rect 2682 22760 2688 22772
rect 2643 22732 2688 22760
rect 2682 22720 2688 22732
rect 2740 22720 2746 22772
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 16758 22760 16764 22772
rect 2832 22732 15700 22760
rect 16719 22732 16764 22760
rect 2832 22720 2838 22732
rect 1670 22652 1676 22704
rect 1728 22692 1734 22704
rect 13078 22692 13084 22704
rect 1728 22664 13084 22692
rect 1728 22652 1734 22664
rect 13078 22652 13084 22664
rect 13136 22652 13142 22704
rect 15672 22692 15700 22732
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 18690 22760 18696 22772
rect 17512 22732 18696 22760
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 15672 22664 17141 22692
rect 17129 22661 17141 22664
rect 17175 22692 17187 22695
rect 17402 22692 17408 22704
rect 17175 22664 17408 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17402 22652 17408 22664
rect 17460 22652 17466 22704
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22624 2651 22627
rect 3510 22624 3516 22636
rect 2639 22596 3516 22624
rect 2639 22593 2651 22596
rect 2593 22587 2651 22593
rect 3510 22584 3516 22596
rect 3568 22584 3574 22636
rect 3970 22633 3976 22636
rect 3964 22587 3976 22633
rect 4028 22624 4034 22636
rect 7098 22624 7104 22636
rect 4028 22596 4064 22624
rect 7059 22596 7104 22624
rect 3970 22584 3976 22587
rect 4028 22584 4034 22596
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 7193 22627 7251 22633
rect 7193 22593 7205 22627
rect 7239 22593 7251 22627
rect 7374 22624 7380 22636
rect 7335 22596 7380 22624
rect 7193 22587 7251 22593
rect 2406 22516 2412 22568
rect 2464 22556 2470 22568
rect 2682 22556 2688 22568
rect 2464 22528 2688 22556
rect 2464 22516 2470 22528
rect 2682 22516 2688 22528
rect 2740 22556 2746 22568
rect 2777 22559 2835 22565
rect 2777 22556 2789 22559
rect 2740 22528 2789 22556
rect 2740 22516 2746 22528
rect 2777 22525 2789 22528
rect 2823 22525 2835 22559
rect 2777 22519 2835 22525
rect 3697 22559 3755 22565
rect 3697 22525 3709 22559
rect 3743 22525 3755 22559
rect 7208 22556 7236 22587
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 11517 22627 11575 22633
rect 7524 22596 7569 22624
rect 7524 22584 7530 22596
rect 11517 22593 11529 22627
rect 11563 22624 11575 22627
rect 14826 22624 14832 22636
rect 11563 22596 14832 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 16942 22624 16948 22636
rect 16903 22596 16948 22624
rect 16942 22584 16948 22596
rect 17000 22584 17006 22636
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22624 17279 22627
rect 17512 22624 17540 22732
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 20346 22760 20352 22772
rect 19352 22732 20352 22760
rect 19352 22692 19380 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 25774 22760 25780 22772
rect 25735 22732 25780 22760
rect 25774 22720 25780 22732
rect 25832 22720 25838 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 25884 22732 26157 22760
rect 18432 22664 19380 22692
rect 18432 22633 18460 22664
rect 24762 22652 24768 22704
rect 24820 22692 24826 22704
rect 25884 22692 25912 22732
rect 26145 22729 26157 22732
rect 26191 22760 26203 22763
rect 26786 22760 26792 22772
rect 26191 22732 26792 22760
rect 26191 22729 26203 22732
rect 26145 22723 26203 22729
rect 26786 22720 26792 22732
rect 26844 22720 26850 22772
rect 27982 22760 27988 22772
rect 27943 22732 27988 22760
rect 27982 22720 27988 22732
rect 28040 22720 28046 22772
rect 32585 22763 32643 22769
rect 32585 22729 32597 22763
rect 32631 22729 32643 22763
rect 32585 22723 32643 22729
rect 26418 22692 26424 22704
rect 24820 22664 25912 22692
rect 25976 22664 26424 22692
rect 24820 22652 24826 22664
rect 17267 22596 17540 22624
rect 18417 22627 18475 22633
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 18509 22627 18567 22633
rect 18509 22593 18521 22627
rect 18555 22624 18567 22627
rect 18966 22624 18972 22636
rect 18555 22596 18972 22624
rect 18555 22593 18567 22596
rect 18509 22587 18567 22593
rect 7742 22556 7748 22568
rect 7208 22528 7748 22556
rect 3697 22519 3755 22525
rect 1486 22448 1492 22500
rect 1544 22488 1550 22500
rect 2314 22488 2320 22500
rect 1544 22460 2320 22488
rect 1544 22448 1550 22460
rect 2314 22448 2320 22460
rect 2372 22488 2378 22500
rect 3712 22488 3740 22519
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 14274 22516 14280 22568
rect 14332 22556 14338 22568
rect 17236 22556 17264 22587
rect 18966 22584 18972 22596
rect 19024 22584 19030 22636
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19518 22624 19524 22636
rect 19208 22596 19380 22624
rect 19479 22596 19524 22624
rect 19208 22584 19214 22596
rect 18598 22556 18604 22568
rect 14332 22528 17264 22556
rect 18559 22528 18604 22556
rect 14332 22516 14338 22528
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 18690 22516 18696 22568
rect 18748 22556 18754 22568
rect 18748 22528 18793 22556
rect 18748 22516 18754 22528
rect 2372 22460 3740 22488
rect 2372 22448 2378 22460
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 5074 22420 5080 22432
rect 5035 22392 5080 22420
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 6917 22423 6975 22429
rect 6917 22389 6929 22423
rect 6963 22420 6975 22423
rect 7006 22420 7012 22432
rect 6963 22392 7012 22420
rect 6963 22389 6975 22392
rect 6917 22383 6975 22389
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 10376 22392 11713 22420
rect 10376 22380 10382 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 13722 22380 13728 22432
rect 13780 22420 13786 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 13780 22392 18245 22420
rect 13780 22380 13786 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 19242 22420 19248 22432
rect 19203 22392 19248 22420
rect 18233 22383 18291 22389
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 19352 22420 19380 22596
rect 19518 22584 19524 22596
rect 19576 22584 19582 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 19794 22624 19800 22636
rect 19751 22596 19800 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 22180 22627 22238 22633
rect 22180 22593 22192 22627
rect 22226 22624 22238 22627
rect 23014 22624 23020 22636
rect 22226 22596 23020 22624
rect 22226 22593 22238 22596
rect 22180 22587 22238 22593
rect 23014 22584 23020 22596
rect 23072 22584 23078 22636
rect 25976 22633 26004 22664
rect 26418 22652 26424 22664
rect 26476 22692 26482 22704
rect 27801 22695 27859 22701
rect 27801 22692 27813 22695
rect 26476 22664 27813 22692
rect 26476 22652 26482 22664
rect 27801 22661 27813 22664
rect 27847 22661 27859 22695
rect 27801 22655 27859 22661
rect 28442 22652 28448 22704
rect 28500 22692 28506 22704
rect 28690 22695 28748 22701
rect 28690 22692 28702 22695
rect 28500 22664 28702 22692
rect 28500 22652 28506 22664
rect 28690 22661 28702 22664
rect 28736 22661 28748 22695
rect 32214 22692 32220 22704
rect 32175 22664 32220 22692
rect 28690 22655 28748 22661
rect 32214 22652 32220 22664
rect 32272 22652 32278 22704
rect 32398 22652 32404 22704
rect 32456 22701 32462 22704
rect 32456 22695 32475 22701
rect 32463 22661 32475 22695
rect 32456 22655 32475 22661
rect 32456 22652 32462 22655
rect 32600 22636 32628 22723
rect 25961 22627 26019 22633
rect 25961 22593 25973 22627
rect 26007 22593 26019 22627
rect 26234 22624 26240 22636
rect 26195 22596 26240 22624
rect 25961 22587 26019 22593
rect 26234 22584 26240 22596
rect 26292 22584 26298 22636
rect 27614 22624 27620 22636
rect 27575 22596 27620 22624
rect 27614 22584 27620 22596
rect 27672 22584 27678 22636
rect 31202 22624 31208 22636
rect 28460 22596 31208 22624
rect 19425 22559 19483 22565
rect 19425 22525 19437 22559
rect 19471 22525 19483 22559
rect 19425 22519 19483 22525
rect 19613 22559 19671 22565
rect 19613 22525 19625 22559
rect 19659 22525 19671 22559
rect 19613 22519 19671 22525
rect 19444 22488 19472 22519
rect 19518 22488 19524 22500
rect 19444 22460 19524 22488
rect 19518 22448 19524 22460
rect 19576 22448 19582 22500
rect 19628 22488 19656 22519
rect 21634 22516 21640 22568
rect 21692 22556 21698 22568
rect 21913 22559 21971 22565
rect 21913 22556 21925 22559
rect 21692 22528 21925 22556
rect 21692 22516 21698 22528
rect 21913 22525 21925 22528
rect 21959 22525 21971 22559
rect 21913 22519 21971 22525
rect 27890 22516 27896 22568
rect 27948 22556 27954 22568
rect 28460 22565 28488 22596
rect 31202 22584 31208 22596
rect 31260 22584 31266 22636
rect 31294 22584 31300 22636
rect 31352 22624 31358 22636
rect 31389 22627 31447 22633
rect 31389 22624 31401 22627
rect 31352 22596 31401 22624
rect 31352 22584 31358 22596
rect 31389 22593 31401 22596
rect 31435 22593 31447 22627
rect 31389 22587 31447 22593
rect 31573 22627 31631 22633
rect 31573 22593 31585 22627
rect 31619 22624 31631 22627
rect 32582 22624 32588 22636
rect 31619 22596 32588 22624
rect 31619 22593 31631 22596
rect 31573 22587 31631 22593
rect 32582 22584 32588 22596
rect 32640 22584 32646 22636
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 33597 22627 33655 22633
rect 33597 22624 33609 22627
rect 33192 22596 33609 22624
rect 33192 22584 33198 22596
rect 33597 22593 33609 22596
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33781 22627 33839 22633
rect 33781 22593 33793 22627
rect 33827 22624 33839 22627
rect 33962 22624 33968 22636
rect 33827 22596 33968 22624
rect 33827 22593 33839 22596
rect 33781 22587 33839 22593
rect 33962 22584 33968 22596
rect 34020 22584 34026 22636
rect 34606 22624 34612 22636
rect 34567 22596 34612 22624
rect 34606 22584 34612 22596
rect 34664 22584 34670 22636
rect 34698 22584 34704 22636
rect 34756 22624 34762 22636
rect 34865 22627 34923 22633
rect 34865 22624 34877 22627
rect 34756 22596 34877 22624
rect 34756 22584 34762 22596
rect 34865 22593 34877 22596
rect 34911 22593 34923 22627
rect 34865 22587 34923 22593
rect 28445 22559 28503 22565
rect 28445 22556 28457 22559
rect 27948 22528 28457 22556
rect 27948 22516 27954 22528
rect 28445 22525 28457 22528
rect 28491 22525 28503 22559
rect 28445 22519 28503 22525
rect 21726 22488 21732 22500
rect 19628 22460 21732 22488
rect 21726 22448 21732 22460
rect 21784 22448 21790 22500
rect 31754 22448 31760 22500
rect 31812 22488 31818 22500
rect 31812 22460 32444 22488
rect 31812 22448 31818 22460
rect 19794 22420 19800 22432
rect 19352 22392 19800 22420
rect 19794 22380 19800 22392
rect 19852 22380 19858 22432
rect 23293 22423 23351 22429
rect 23293 22389 23305 22423
rect 23339 22420 23351 22423
rect 23382 22420 23388 22432
rect 23339 22392 23388 22420
rect 23339 22389 23351 22392
rect 23293 22383 23351 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 29825 22423 29883 22429
rect 29825 22389 29837 22423
rect 29871 22420 29883 22423
rect 30190 22420 30196 22432
rect 29871 22392 30196 22420
rect 29871 22389 29883 22392
rect 29825 22383 29883 22389
rect 30190 22380 30196 22392
rect 30248 22380 30254 22432
rect 31389 22423 31447 22429
rect 31389 22389 31401 22423
rect 31435 22420 31447 22423
rect 31938 22420 31944 22432
rect 31435 22392 31944 22420
rect 31435 22389 31447 22392
rect 31389 22383 31447 22389
rect 31938 22380 31944 22392
rect 31996 22380 32002 22432
rect 32416 22429 32444 22460
rect 32401 22423 32459 22429
rect 32401 22389 32413 22423
rect 32447 22420 32459 22423
rect 32766 22420 32772 22432
rect 32447 22392 32772 22420
rect 32447 22389 32459 22392
rect 32401 22383 32459 22389
rect 32766 22380 32772 22392
rect 32824 22380 32830 22432
rect 33965 22423 34023 22429
rect 33965 22389 33977 22423
rect 34011 22420 34023 22423
rect 34790 22420 34796 22432
rect 34011 22392 34796 22420
rect 34011 22389 34023 22392
rect 33965 22383 34023 22389
rect 34790 22380 34796 22392
rect 34848 22380 34854 22432
rect 35989 22423 36047 22429
rect 35989 22389 36001 22423
rect 36035 22420 36047 22423
rect 36262 22420 36268 22432
rect 36035 22392 36268 22420
rect 36035 22389 36047 22392
rect 35989 22383 36047 22389
rect 36262 22380 36268 22392
rect 36320 22380 36326 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1394 22176 1400 22228
rect 1452 22216 1458 22228
rect 11977 22219 12035 22225
rect 11977 22216 11989 22219
rect 1452 22188 11989 22216
rect 1452 22176 1458 22188
rect 11977 22185 11989 22188
rect 12023 22185 12035 22219
rect 19242 22216 19248 22228
rect 11977 22179 12035 22185
rect 18340 22188 19248 22216
rect 2682 22108 2688 22160
rect 2740 22148 2746 22160
rect 2740 22120 4476 22148
rect 2740 22108 2746 22120
rect 4448 22094 4476 22120
rect 4448 22089 4513 22094
rect 4433 22083 4513 22089
rect 4433 22049 4445 22083
rect 4479 22066 4513 22083
rect 4479 22049 4491 22066
rect 4433 22043 4491 22049
rect 7098 22040 7104 22092
rect 7156 22080 7162 22092
rect 7156 22052 7512 22080
rect 7156 22040 7162 22052
rect 1854 22012 1860 22024
rect 1815 21984 1860 22012
rect 1854 21972 1860 21984
rect 1912 21972 1918 22024
rect 2866 22012 2872 22024
rect 2827 21984 2872 22012
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 5074 22012 5080 22024
rect 4295 21984 5080 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 6696 21984 7205 22012
rect 6696 21972 6702 21984
rect 7193 21981 7205 21984
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 7484 22021 7512 22052
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 10226 22080 10232 22092
rect 9732 22052 10232 22080
rect 9732 22040 9738 22052
rect 10226 22040 10232 22052
rect 10284 22080 10290 22092
rect 10597 22083 10655 22089
rect 10597 22080 10609 22083
rect 10284 22052 10609 22080
rect 10284 22040 10290 22052
rect 10597 22049 10609 22052
rect 10643 22049 10655 22083
rect 11992 22080 12020 22179
rect 11992 22052 12848 22080
rect 10597 22043 10655 22049
rect 12820 22021 12848 22052
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 13044 22052 14105 22080
rect 13044 22040 13050 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 18141 22083 18199 22089
rect 18141 22049 18153 22083
rect 18187 22080 18199 22083
rect 18230 22080 18236 22092
rect 18187 22052 18236 22080
rect 18187 22049 18199 22052
rect 18141 22043 18199 22049
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 18340 22089 18368 22188
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 20346 22216 20352 22228
rect 20307 22188 20352 22216
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 20806 22216 20812 22228
rect 20456 22188 20812 22216
rect 18598 22148 18604 22160
rect 18524 22120 18604 22148
rect 18524 22089 18552 22120
rect 18598 22108 18604 22120
rect 18656 22108 18662 22160
rect 18874 22108 18880 22160
rect 18932 22148 18938 22160
rect 19337 22151 19395 22157
rect 19337 22148 19349 22151
rect 18932 22120 19349 22148
rect 18932 22108 18938 22120
rect 19337 22117 19349 22120
rect 19383 22117 19395 22151
rect 19978 22148 19984 22160
rect 19337 22111 19395 22117
rect 19629 22120 19984 22148
rect 18325 22083 18383 22089
rect 18325 22049 18337 22083
rect 18371 22049 18383 22083
rect 18325 22043 18383 22049
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22080 18567 22083
rect 18555 22052 18589 22080
rect 18555 22049 18567 22052
rect 18509 22043 18567 22049
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19629 22080 19657 22120
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 19576 22052 19669 22080
rect 19576 22040 19582 22052
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 20456 22080 20484 22188
rect 20806 22176 20812 22188
rect 20864 22176 20870 22228
rect 23014 22216 23020 22228
rect 22975 22188 23020 22216
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 27614 22176 27620 22228
rect 27672 22216 27678 22228
rect 28353 22219 28411 22225
rect 28353 22216 28365 22219
rect 27672 22188 28365 22216
rect 27672 22176 27678 22188
rect 28353 22185 28365 22188
rect 28399 22185 28411 22219
rect 28353 22179 28411 22185
rect 28442 22176 28448 22228
rect 28500 22216 28506 22228
rect 31478 22216 31484 22228
rect 28500 22188 29040 22216
rect 31439 22188 31484 22216
rect 28500 22176 28506 22188
rect 23382 22148 23388 22160
rect 20732 22120 23388 22148
rect 20622 22080 20628 22092
rect 19852 22052 20484 22080
rect 20583 22052 20628 22080
rect 19852 22040 19858 22052
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 20732 22089 20760 22120
rect 23382 22108 23388 22120
rect 23440 22108 23446 22160
rect 28810 22108 28816 22160
rect 28868 22108 28874 22160
rect 28902 22108 28908 22160
rect 28960 22108 28966 22160
rect 20717 22083 20775 22089
rect 20717 22049 20729 22083
rect 20763 22049 20775 22083
rect 28828 22080 28856 22108
rect 20717 22043 20775 22049
rect 28736 22052 28856 22080
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 7929 22015 7987 22021
rect 7929 21981 7941 22015
rect 7975 21981 7987 22015
rect 7929 21975 7987 21981
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 2225 21947 2283 21953
rect 2225 21913 2237 21947
rect 2271 21944 2283 21947
rect 2314 21944 2320 21956
rect 2271 21916 2320 21944
rect 2271 21913 2283 21916
rect 2225 21907 2283 21913
rect 2314 21904 2320 21916
rect 2372 21904 2378 21956
rect 4341 21947 4399 21953
rect 4341 21944 4353 21947
rect 2700 21916 4353 21944
rect 2700 21885 2728 21916
rect 4341 21913 4353 21916
rect 4387 21913 4399 21947
rect 4341 21907 4399 21913
rect 7098 21904 7104 21956
rect 7156 21944 7162 21956
rect 7392 21944 7420 21972
rect 7944 21944 7972 21975
rect 8202 21944 8208 21956
rect 7156 21916 7420 21944
rect 7484 21916 8208 21944
rect 7156 21904 7162 21916
rect 7484 21888 7512 21916
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 10864 21947 10922 21953
rect 10864 21913 10876 21947
rect 10910 21944 10922 21947
rect 12437 21947 12495 21953
rect 12437 21944 12449 21947
rect 10910 21916 12449 21944
rect 10910 21913 10922 21916
rect 10864 21907 10922 21913
rect 12437 21913 12449 21916
rect 12483 21913 12495 21947
rect 12437 21907 12495 21913
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21845 2743 21879
rect 3878 21876 3884 21888
rect 3839 21848 3884 21876
rect 2685 21839 2743 21845
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 7006 21876 7012 21888
rect 6967 21848 7012 21876
rect 7006 21836 7012 21848
rect 7064 21836 7070 21888
rect 7377 21879 7435 21885
rect 7377 21845 7389 21879
rect 7423 21876 7435 21879
rect 7466 21876 7472 21888
rect 7423 21848 7472 21876
rect 7423 21845 7435 21848
rect 7377 21839 7435 21845
rect 7466 21836 7472 21848
rect 7524 21836 7530 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 8113 21879 8171 21885
rect 8113 21876 8125 21879
rect 7800 21848 8125 21876
rect 7800 21836 7806 21848
rect 8113 21845 8125 21848
rect 8159 21845 8171 21879
rect 12636 21876 12664 21975
rect 12894 21972 12900 22024
rect 12952 22012 12958 22024
rect 14182 22012 14188 22024
rect 12952 21984 14188 22012
rect 12952 21972 12958 21984
rect 14182 21972 14188 21984
rect 14240 21972 14246 22024
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 18601 22015 18659 22021
rect 18601 21981 18613 22015
rect 18647 22012 18659 22015
rect 18690 22012 18696 22024
rect 18647 21984 18696 22012
rect 18647 21981 18659 21984
rect 18601 21975 18659 21981
rect 13814 21904 13820 21956
rect 13872 21944 13878 21956
rect 14338 21947 14396 21953
rect 14338 21944 14350 21947
rect 13872 21916 14350 21944
rect 13872 21904 13878 21916
rect 14338 21913 14350 21916
rect 14384 21913 14396 21947
rect 18432 21944 18460 21975
rect 18690 21972 18696 21984
rect 18748 21972 18754 22024
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 19426 22012 19432 22024
rect 18840 21984 19432 22012
rect 18840 21972 18846 21984
rect 19426 21972 19432 21984
rect 19484 22012 19490 22024
rect 19613 22015 19671 22021
rect 19613 22012 19625 22015
rect 19484 21984 19625 22012
rect 19484 21972 19490 21984
rect 19613 21981 19625 21984
rect 19659 21981 19671 22015
rect 19613 21975 19671 21981
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20438 22012 20444 22024
rect 19751 21984 20444 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20806 22012 20812 22024
rect 20579 21984 20668 22012
rect 20767 21984 20812 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20346 21944 20352 21956
rect 18432 21916 20352 21944
rect 14338 21907 14396 21913
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 15194 21876 15200 21888
rect 12636 21848 15200 21876
rect 8113 21839 8171 21845
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 15470 21876 15476 21888
rect 15431 21848 15476 21876
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 20640 21876 20668 21984
rect 20806 21972 20812 21984
rect 20864 21972 20870 22024
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22370 22012 22376 22024
rect 22327 21984 22376 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22520 21984 22569 22012
rect 22520 21972 22526 21984
rect 22557 21981 22569 21984
rect 22603 22012 22615 22015
rect 23106 22012 23112 22024
rect 22603 21984 23112 22012
rect 22603 21981 22615 21984
rect 22557 21975 22615 21981
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 22012 23259 22015
rect 23477 22015 23535 22021
rect 23247 21981 23263 22012
rect 23201 21975 23263 21981
rect 23477 21981 23489 22015
rect 23523 22012 23535 22015
rect 26234 22012 26240 22024
rect 23523 21984 26240 22012
rect 23523 21981 23535 21984
rect 23477 21975 23535 21981
rect 21726 21904 21732 21956
rect 21784 21944 21790 21956
rect 23235 21944 23263 21975
rect 23382 21944 23388 21956
rect 21784 21916 22508 21944
rect 21784 21904 21790 21916
rect 17920 21848 20668 21876
rect 17920 21836 17926 21848
rect 22094 21836 22100 21888
rect 22152 21876 22158 21888
rect 22480 21885 22508 21916
rect 23216 21916 23263 21944
rect 23343 21916 23388 21944
rect 22465 21879 22523 21885
rect 22152 21848 22197 21876
rect 22152 21836 22158 21848
rect 22465 21845 22477 21879
rect 22511 21845 22523 21879
rect 22465 21839 22523 21845
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 23216 21876 23244 21916
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 23072 21848 23244 21876
rect 23072 21836 23078 21848
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 23492 21876 23520 21975
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 28736 22021 28764 22052
rect 28629 22015 28687 22021
rect 28629 21981 28641 22015
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 28721 22015 28779 22021
rect 28721 21981 28733 22015
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 22012 28871 22015
rect 28920 22012 28948 22108
rect 29012 22080 29040 22188
rect 31478 22176 31484 22188
rect 31536 22176 31542 22228
rect 34698 22216 34704 22228
rect 34659 22188 34704 22216
rect 34698 22176 34704 22188
rect 34756 22176 34762 22228
rect 30190 22108 30196 22160
rect 30248 22148 30254 22160
rect 32030 22148 32036 22160
rect 30248 22120 32036 22148
rect 30248 22108 30254 22120
rect 32030 22108 32036 22120
rect 32088 22108 32094 22160
rect 32953 22083 33011 22089
rect 29012 22052 32536 22080
rect 28859 21984 28948 22012
rect 28997 22015 29055 22021
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 28997 21981 29009 22015
rect 29043 22012 29055 22015
rect 29086 22012 29092 22024
rect 29043 21984 29092 22012
rect 29043 21981 29055 21984
rect 28997 21975 29055 21981
rect 28644 21944 28672 21975
rect 29086 21972 29092 21984
rect 29144 21972 29150 22024
rect 30190 22012 30196 22024
rect 30151 21984 30196 22012
rect 30190 21972 30196 21984
rect 30248 21972 30254 22024
rect 30469 22015 30527 22021
rect 30469 21981 30481 22015
rect 30515 21981 30527 22015
rect 30469 21975 30527 21981
rect 29178 21944 29184 21956
rect 28644 21916 29184 21944
rect 29178 21904 29184 21916
rect 29236 21944 29242 21956
rect 30484 21944 30512 21975
rect 30558 21972 30564 22024
rect 30616 22012 30622 22024
rect 31386 22012 31392 22024
rect 30616 21984 31392 22012
rect 30616 21972 30622 21984
rect 31386 21972 31392 21984
rect 31444 22012 31450 22024
rect 31665 22015 31723 22021
rect 31665 22012 31677 22015
rect 31444 21984 31677 22012
rect 31444 21972 31450 21984
rect 31665 21981 31677 21984
rect 31711 21981 31723 22015
rect 31938 22012 31944 22024
rect 31899 21984 31944 22012
rect 31665 21975 31723 21981
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 31478 21944 31484 21956
rect 29236 21916 31484 21944
rect 29236 21904 29242 21916
rect 31478 21904 31484 21916
rect 31536 21904 31542 21956
rect 31846 21876 31852 21888
rect 23348 21848 23520 21876
rect 31807 21848 31852 21876
rect 23348 21836 23354 21848
rect 31846 21836 31852 21848
rect 31904 21836 31910 21888
rect 32508 21876 32536 22052
rect 32953 22049 32965 22083
rect 32999 22080 33011 22083
rect 33134 22080 33140 22092
rect 32999 22052 33140 22080
rect 32999 22049 33011 22052
rect 32953 22043 33011 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 36262 22080 36268 22092
rect 33244 22052 36268 22080
rect 32674 21972 32680 22024
rect 32732 22012 32738 22024
rect 33244 22021 33272 22052
rect 36262 22040 36268 22052
rect 36320 22040 36326 22092
rect 33229 22015 33287 22021
rect 33229 22012 33241 22015
rect 32732 21984 33241 22012
rect 32732 21972 32738 21984
rect 33229 21981 33241 21984
rect 33275 21981 33287 22015
rect 33229 21975 33287 21981
rect 33321 22015 33379 22021
rect 33321 21981 33333 22015
rect 33367 21981 33379 22015
rect 33321 21975 33379 21981
rect 32582 21904 32588 21956
rect 32640 21944 32646 21956
rect 33336 21944 33364 21975
rect 33410 21972 33416 22024
rect 33468 22012 33474 22024
rect 33468 21984 33513 22012
rect 33468 21972 33474 21984
rect 33594 21972 33600 22024
rect 33652 22012 33658 22024
rect 33652 21984 33697 22012
rect 33652 21972 33658 21984
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34848 21984 34897 22012
rect 34848 21972 34854 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 37921 22015 37979 22021
rect 37921 21981 37933 22015
rect 37967 22012 37979 22015
rect 39114 22012 39120 22024
rect 37967 21984 39120 22012
rect 37967 21981 37979 21984
rect 37921 21975 37979 21981
rect 39114 21972 39120 21984
rect 39172 21972 39178 22024
rect 32640 21916 33364 21944
rect 32640 21904 32646 21916
rect 34422 21904 34428 21956
rect 34480 21944 34486 21956
rect 37826 21944 37832 21956
rect 34480 21916 37832 21944
rect 34480 21904 34486 21916
rect 37826 21904 37832 21916
rect 37884 21904 37890 21956
rect 38188 21947 38246 21953
rect 38188 21913 38200 21947
rect 38234 21944 38246 21947
rect 38286 21944 38292 21956
rect 38234 21916 38292 21944
rect 38234 21913 38246 21916
rect 38188 21907 38246 21913
rect 38286 21904 38292 21916
rect 38344 21904 38350 21956
rect 35710 21876 35716 21888
rect 32508 21848 35716 21876
rect 35710 21836 35716 21848
rect 35768 21836 35774 21888
rect 38654 21836 38660 21888
rect 38712 21876 38718 21888
rect 39301 21879 39359 21885
rect 39301 21876 39313 21879
rect 38712 21848 39313 21876
rect 38712 21836 38718 21848
rect 39301 21845 39313 21848
rect 39347 21845 39359 21879
rect 39301 21839 39359 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 3881 21675 3939 21681
rect 3881 21641 3893 21675
rect 3927 21672 3939 21675
rect 3970 21672 3976 21684
rect 3927 21644 3976 21672
rect 3927 21641 3939 21644
rect 3881 21635 3939 21641
rect 3970 21632 3976 21644
rect 4028 21632 4034 21684
rect 7098 21632 7104 21684
rect 7156 21672 7162 21684
rect 7282 21672 7288 21684
rect 7156 21644 7288 21672
rect 7156 21632 7162 21644
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 7558 21632 7564 21684
rect 7616 21672 7622 21684
rect 7742 21672 7748 21684
rect 7616 21644 7748 21672
rect 7616 21632 7622 21644
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 13814 21672 13820 21684
rect 13775 21644 13820 21672
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 16632 21644 16681 21672
rect 16632 21632 16638 21644
rect 16669 21641 16681 21644
rect 16715 21641 16727 21675
rect 16669 21635 16727 21641
rect 18414 21632 18420 21684
rect 18472 21672 18478 21684
rect 19061 21675 19119 21681
rect 19061 21672 19073 21675
rect 18472 21644 19073 21672
rect 18472 21632 18478 21644
rect 19061 21641 19073 21644
rect 19107 21641 19119 21675
rect 19061 21635 19119 21641
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 24762 21672 24768 21684
rect 20496 21644 24768 21672
rect 20496 21632 20502 21644
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 28902 21632 28908 21684
rect 28960 21672 28966 21684
rect 29089 21675 29147 21681
rect 29089 21672 29101 21675
rect 28960 21644 29101 21672
rect 28960 21632 28966 21644
rect 29089 21641 29101 21644
rect 29135 21641 29147 21675
rect 30558 21672 30564 21684
rect 29089 21635 29147 21641
rect 29196 21644 30564 21672
rect 14185 21607 14243 21613
rect 14185 21604 14197 21607
rect 1412 21576 14197 21604
rect 1412 21545 1440 21576
rect 14185 21573 14197 21576
rect 14231 21604 14243 21607
rect 15470 21604 15476 21616
rect 14231 21576 15476 21604
rect 14231 21573 14243 21576
rect 14185 21567 14243 21573
rect 15470 21564 15476 21576
rect 15528 21564 15534 21616
rect 15562 21564 15568 21616
rect 15620 21604 15626 21616
rect 15620 21576 18552 21604
rect 15620 21564 15626 21576
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 2038 21536 2044 21548
rect 1820 21508 2044 21536
rect 1820 21496 1826 21508
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 2406 21536 2412 21548
rect 2367 21508 2412 21536
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 3050 21536 3056 21548
rect 3011 21508 3056 21536
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 3878 21496 3884 21548
rect 3936 21536 3942 21548
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 3936 21508 4077 21536
rect 3936 21496 3942 21508
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21505 6975 21539
rect 7190 21536 7196 21548
rect 7151 21508 7196 21536
rect 6917 21499 6975 21505
rect 6932 21400 6960 21499
rect 7190 21496 7196 21508
rect 7248 21496 7254 21548
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7742 21536 7748 21548
rect 7340 21508 7748 21536
rect 7340 21496 7346 21508
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21536 7895 21539
rect 8110 21536 8116 21548
rect 7883 21508 8116 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 8110 21496 8116 21508
rect 8168 21496 8174 21548
rect 8202 21496 8208 21548
rect 8260 21536 8266 21548
rect 8665 21539 8723 21545
rect 8665 21536 8677 21539
rect 8260 21508 8677 21536
rect 8260 21496 8266 21508
rect 8665 21505 8677 21508
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 14001 21539 14059 21545
rect 14001 21505 14013 21539
rect 14047 21505 14059 21539
rect 14274 21536 14280 21548
rect 14235 21508 14280 21536
rect 14001 21499 14059 21505
rect 7098 21468 7104 21480
rect 7059 21440 7104 21468
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 7208 21468 7236 21496
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7208 21440 7941 21468
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 8018 21428 8024 21480
rect 8076 21468 8082 21480
rect 8864 21468 8892 21499
rect 8076 21440 8892 21468
rect 8076 21428 8082 21440
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 6932 21372 8769 21400
rect 8757 21369 8769 21372
rect 8803 21369 8815 21403
rect 8757 21363 8815 21369
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 2222 21332 2228 21344
rect 2183 21304 2228 21332
rect 2222 21292 2228 21304
rect 2280 21292 2286 21344
rect 2866 21332 2872 21344
rect 2827 21304 2872 21332
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7193 21335 7251 21341
rect 7193 21332 7205 21335
rect 6972 21304 7205 21332
rect 6972 21292 6978 21304
rect 7193 21301 7205 21304
rect 7239 21332 7251 21335
rect 7282 21332 7288 21344
rect 7239 21304 7288 21332
rect 7239 21301 7251 21304
rect 7193 21295 7251 21301
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7377 21335 7435 21341
rect 7377 21301 7389 21335
rect 7423 21332 7435 21335
rect 7742 21332 7748 21344
rect 7423 21304 7748 21332
rect 7423 21301 7435 21304
rect 7377 21295 7435 21301
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 8202 21332 8208 21344
rect 7892 21304 7937 21332
rect 8163 21304 8208 21332
rect 7892 21292 7898 21304
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 14016 21332 14044 21499
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 14608 21508 14841 21536
rect 14608 21496 14614 21508
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 14829 21499 14887 21505
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16632 21508 17049 21536
rect 16632 21496 16638 21508
rect 17037 21505 17049 21508
rect 17083 21536 17095 21539
rect 17586 21536 17592 21548
rect 17083 21508 17592 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 17954 21536 17960 21548
rect 17915 21508 17960 21536
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 18524 21536 18552 21576
rect 18598 21564 18604 21616
rect 18656 21604 18662 21616
rect 18656 21576 19472 21604
rect 18656 21564 18662 21576
rect 18782 21536 18788 21548
rect 18524 21508 18788 21536
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 18874 21496 18880 21548
rect 18932 21536 18938 21548
rect 19444 21545 19472 21576
rect 22370 21564 22376 21616
rect 22428 21604 22434 21616
rect 29196 21604 29224 21644
rect 30558 21632 30564 21644
rect 30616 21632 30622 21684
rect 31478 21672 31484 21684
rect 31439 21644 31484 21672
rect 31478 21632 31484 21644
rect 31536 21632 31542 21684
rect 31570 21632 31576 21684
rect 31628 21672 31634 21684
rect 33045 21675 33103 21681
rect 33045 21672 33057 21675
rect 31628 21644 33057 21672
rect 31628 21632 31634 21644
rect 33045 21641 33057 21644
rect 33091 21641 33103 21675
rect 33045 21635 33103 21641
rect 33410 21632 33416 21684
rect 33468 21672 33474 21684
rect 33781 21675 33839 21681
rect 33781 21672 33793 21675
rect 33468 21644 33793 21672
rect 33468 21632 33474 21644
rect 33781 21641 33793 21644
rect 33827 21641 33839 21675
rect 35710 21672 35716 21684
rect 35671 21644 35716 21672
rect 33781 21635 33839 21641
rect 35710 21632 35716 21644
rect 35768 21632 35774 21684
rect 22428 21576 29224 21604
rect 22428 21564 22434 21576
rect 32030 21564 32036 21616
rect 32088 21604 32094 21616
rect 32953 21607 33011 21613
rect 32953 21604 32965 21607
rect 32088 21576 32965 21604
rect 32088 21564 32094 21576
rect 32953 21573 32965 21576
rect 32999 21573 33011 21607
rect 32953 21567 33011 21573
rect 35250 21564 35256 21616
rect 35308 21604 35314 21616
rect 35345 21607 35403 21613
rect 35345 21604 35357 21607
rect 35308 21576 35357 21604
rect 35308 21564 35314 21576
rect 35345 21573 35357 21576
rect 35391 21573 35403 21607
rect 35345 21567 35403 21573
rect 35802 21564 35808 21616
rect 35860 21604 35866 21616
rect 36265 21607 36323 21613
rect 36265 21604 36277 21607
rect 35860 21576 36277 21604
rect 35860 21564 35866 21576
rect 36265 21573 36277 21576
rect 36311 21573 36323 21607
rect 36265 21567 36323 21573
rect 19245 21539 19303 21545
rect 19245 21536 19257 21539
rect 18932 21508 19257 21536
rect 18932 21496 18938 21508
rect 19245 21505 19257 21508
rect 19291 21505 19303 21539
rect 19245 21499 19303 21505
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 24940 21539 24998 21545
rect 24940 21505 24952 21539
rect 24986 21536 24998 21539
rect 25222 21536 25228 21548
rect 24986 21508 25228 21536
rect 24986 21505 24998 21508
rect 24940 21499 24998 21505
rect 25222 21496 25228 21508
rect 25280 21496 25286 21548
rect 28810 21496 28816 21548
rect 28868 21536 28874 21548
rect 28997 21539 29055 21545
rect 28997 21536 29009 21539
rect 28868 21508 29009 21536
rect 28868 21496 28874 21508
rect 28997 21505 29009 21508
rect 29043 21505 29055 21539
rect 29178 21536 29184 21548
rect 29139 21508 29184 21536
rect 28997 21499 29055 21505
rect 29178 21496 29184 21508
rect 29236 21496 29242 21548
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31588 21545 31754 21546
rect 31297 21539 31355 21545
rect 31573 21542 31754 21545
rect 31297 21536 31309 21539
rect 31168 21508 31309 21536
rect 31168 21496 31174 21508
rect 31297 21505 31309 21508
rect 31343 21505 31355 21539
rect 31487 21539 31754 21542
rect 31487 21536 31585 21539
rect 31297 21499 31355 21505
rect 31404 21514 31585 21536
rect 31404 21508 31515 21514
rect 15654 21428 15660 21480
rect 15712 21468 15718 21480
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 15712 21440 16865 21468
rect 15712 21428 15718 21440
rect 16853 21437 16865 21440
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17129 21471 17187 21477
rect 17000 21440 17045 21468
rect 17000 21428 17006 21440
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 17678 21468 17684 21480
rect 17175 21440 17684 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 17862 21468 17868 21480
rect 17823 21440 17868 21468
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21437 18107 21471
rect 18049 21431 18107 21437
rect 15013 21403 15071 21409
rect 15013 21369 15025 21403
rect 15059 21400 15071 21403
rect 15838 21400 15844 21412
rect 15059 21372 15844 21400
rect 15059 21369 15071 21372
rect 15013 21363 15071 21369
rect 15838 21360 15844 21372
rect 15896 21360 15902 21412
rect 18064 21400 18092 21431
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 19150 21468 19156 21480
rect 18196 21440 19156 21468
rect 18196 21428 18202 21440
rect 19150 21428 19156 21440
rect 19208 21428 19214 21480
rect 19334 21468 19340 21480
rect 19295 21440 19340 21468
rect 19334 21428 19340 21440
rect 19392 21428 19398 21480
rect 19521 21471 19579 21477
rect 19521 21437 19533 21471
rect 19567 21468 19579 21471
rect 20070 21468 20076 21480
rect 19567 21440 20076 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 24394 21428 24400 21480
rect 24452 21468 24458 21480
rect 24670 21468 24676 21480
rect 24452 21440 24676 21468
rect 24452 21428 24458 21440
rect 24670 21428 24676 21440
rect 24728 21428 24734 21480
rect 31404 21468 31432 21508
rect 31573 21505 31585 21514
rect 31619 21518 31754 21539
rect 32674 21536 32680 21548
rect 31619 21505 31631 21518
rect 31573 21499 31631 21505
rect 28966 21440 31432 21468
rect 31726 21468 31754 21518
rect 32635 21508 32680 21536
rect 32674 21496 32680 21508
rect 32732 21496 32738 21548
rect 32858 21496 32864 21548
rect 32916 21536 32922 21548
rect 33229 21539 33287 21545
rect 32916 21508 33009 21536
rect 32916 21496 32922 21508
rect 33229 21505 33241 21539
rect 33275 21536 33287 21539
rect 33686 21536 33692 21548
rect 33275 21508 33692 21536
rect 33275 21505 33287 21508
rect 33229 21499 33287 21505
rect 33686 21496 33692 21508
rect 33744 21496 33750 21548
rect 34698 21496 34704 21548
rect 34756 21536 34762 21548
rect 34880 21545 35112 21546
rect 34880 21539 35127 21545
rect 34880 21536 35081 21539
rect 34756 21518 35081 21536
rect 34756 21508 34908 21518
rect 34756 21496 34762 21508
rect 35069 21505 35081 21518
rect 35115 21505 35127 21539
rect 35069 21499 35127 21505
rect 35162 21539 35220 21545
rect 35162 21505 35174 21539
rect 35208 21505 35220 21539
rect 35162 21499 35220 21505
rect 32398 21468 32404 21480
rect 31726 21440 32404 21468
rect 22370 21400 22376 21412
rect 18064 21372 22376 21400
rect 22370 21360 22376 21372
rect 22428 21360 22434 21412
rect 16206 21332 16212 21344
rect 14016 21304 16212 21332
rect 16206 21292 16212 21304
rect 16264 21292 16270 21344
rect 17402 21292 17408 21344
rect 17460 21332 17466 21344
rect 17681 21335 17739 21341
rect 17681 21332 17693 21335
rect 17460 21304 17693 21332
rect 17460 21292 17466 21304
rect 17681 21301 17693 21304
rect 17727 21301 17739 21335
rect 17681 21295 17739 21301
rect 18966 21292 18972 21344
rect 19024 21332 19030 21344
rect 25958 21332 25964 21344
rect 19024 21304 25964 21332
rect 19024 21292 19030 21304
rect 25958 21292 25964 21304
rect 26016 21292 26022 21344
rect 26050 21292 26056 21344
rect 26108 21332 26114 21344
rect 26108 21304 26153 21332
rect 26108 21292 26114 21304
rect 27246 21292 27252 21344
rect 27304 21332 27310 21344
rect 28258 21332 28264 21344
rect 27304 21304 28264 21332
rect 27304 21292 27310 21304
rect 28258 21292 28264 21304
rect 28316 21292 28322 21344
rect 28810 21292 28816 21344
rect 28868 21332 28874 21344
rect 28966 21332 28994 21440
rect 32398 21428 32404 21440
rect 32456 21468 32462 21480
rect 32582 21468 32588 21480
rect 32456 21440 32588 21468
rect 32456 21428 32462 21440
rect 32582 21428 32588 21440
rect 32640 21428 32646 21480
rect 32876 21468 32904 21496
rect 35177 21468 35205 21499
rect 35434 21496 35440 21548
rect 35492 21536 35498 21548
rect 35575 21539 35633 21545
rect 35492 21508 35537 21536
rect 35492 21496 35498 21508
rect 35575 21505 35587 21539
rect 35621 21536 35633 21539
rect 36170 21536 36176 21548
rect 35621 21508 36176 21536
rect 35621 21505 35633 21508
rect 35575 21499 35633 21505
rect 36170 21496 36176 21508
rect 36228 21496 36234 21548
rect 38654 21496 38660 21548
rect 38712 21536 38718 21548
rect 38749 21539 38807 21545
rect 38749 21536 38761 21539
rect 38712 21508 38761 21536
rect 38712 21496 38718 21508
rect 38749 21505 38761 21508
rect 38795 21505 38807 21539
rect 38749 21499 38807 21505
rect 38838 21468 38844 21480
rect 32876 21440 35205 21468
rect 38799 21440 38844 21468
rect 38838 21428 38844 21440
rect 38896 21428 38902 21480
rect 31294 21400 31300 21412
rect 31255 21372 31300 21400
rect 31294 21360 31300 21372
rect 31352 21360 31358 21412
rect 34790 21360 34796 21412
rect 34848 21400 34854 21412
rect 35526 21400 35532 21412
rect 34848 21372 35532 21400
rect 34848 21360 34854 21372
rect 35526 21360 35532 21372
rect 35584 21400 35590 21412
rect 35802 21400 35808 21412
rect 35584 21372 35808 21400
rect 35584 21360 35590 21372
rect 35802 21360 35808 21372
rect 35860 21360 35866 21412
rect 36449 21403 36507 21409
rect 36449 21369 36461 21403
rect 36495 21400 36507 21403
rect 38010 21400 38016 21412
rect 36495 21372 38016 21400
rect 36495 21369 36507 21372
rect 36449 21363 36507 21369
rect 38010 21360 38016 21372
rect 38068 21360 38074 21412
rect 28868 21304 28994 21332
rect 28868 21292 28874 21304
rect 31846 21292 31852 21344
rect 31904 21332 31910 21344
rect 33410 21332 33416 21344
rect 31904 21304 33416 21332
rect 31904 21292 31910 21304
rect 33410 21292 33416 21304
rect 33468 21332 33474 21344
rect 34422 21332 34428 21344
rect 33468 21304 34428 21332
rect 33468 21292 33474 21304
rect 34422 21292 34428 21304
rect 34480 21292 34486 21344
rect 34606 21292 34612 21344
rect 34664 21332 34670 21344
rect 35434 21332 35440 21344
rect 34664 21304 35440 21332
rect 34664 21292 34670 21304
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 38746 21292 38752 21344
rect 38804 21332 38810 21344
rect 39025 21335 39083 21341
rect 39025 21332 39037 21335
rect 38804 21304 39037 21332
rect 38804 21292 38810 21304
rect 39025 21301 39037 21304
rect 39071 21301 39083 21335
rect 39025 21295 39083 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 7742 21128 7748 21140
rect 7703 21100 7748 21128
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 7834 21088 7840 21140
rect 7892 21128 7898 21140
rect 14550 21128 14556 21140
rect 7892 21100 14556 21128
rect 7892 21088 7898 21100
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 15654 21128 15660 21140
rect 15615 21100 15660 21128
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 16850 21088 16856 21140
rect 16908 21128 16914 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 16908 21100 17233 21128
rect 16908 21088 16914 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 17586 21088 17592 21140
rect 17644 21128 17650 21140
rect 18598 21128 18604 21140
rect 17644 21100 18604 21128
rect 17644 21088 17650 21100
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 25222 21128 25228 21140
rect 19392 21100 25084 21128
rect 25183 21100 25228 21128
rect 19392 21088 19398 21100
rect 7561 21063 7619 21069
rect 7561 21029 7573 21063
rect 7607 21060 7619 21063
rect 7650 21060 7656 21072
rect 7607 21032 7656 21060
rect 7607 21029 7619 21032
rect 7561 21023 7619 21029
rect 7650 21020 7656 21032
rect 7708 21020 7714 21072
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 19245 21063 19303 21069
rect 19245 21060 19257 21063
rect 9364 21032 19257 21060
rect 9364 21020 9370 21032
rect 19245 21029 19257 21032
rect 19291 21029 19303 21063
rect 19610 21060 19616 21072
rect 19245 21023 19303 21029
rect 19352 21032 19616 21060
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 1673 20995 1731 21001
rect 1673 20992 1685 20995
rect 1544 20964 1685 20992
rect 1544 20952 1550 20964
rect 1673 20961 1685 20964
rect 1719 20961 1731 20995
rect 1673 20955 1731 20961
rect 2866 20952 2872 21004
rect 2924 20992 2930 21004
rect 13354 20992 13360 21004
rect 2924 20964 13360 20992
rect 2924 20952 2930 20964
rect 13354 20952 13360 20964
rect 13412 20952 13418 21004
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 15712 20964 15945 20992
rect 15712 20952 15718 20964
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 17402 20992 17408 21004
rect 17363 20964 17408 20992
rect 15933 20955 15991 20961
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17586 20992 17592 21004
rect 17547 20964 17592 20992
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 19352 20992 19380 21032
rect 19610 21020 19616 21032
rect 19668 21020 19674 21072
rect 25056 21060 25084 21100
rect 25222 21088 25228 21100
rect 25280 21088 25286 21140
rect 25958 21088 25964 21140
rect 26016 21128 26022 21140
rect 36817 21131 36875 21137
rect 36817 21128 36829 21131
rect 26016 21100 36829 21128
rect 26016 21088 26022 21100
rect 36817 21097 36829 21100
rect 36863 21097 36875 21131
rect 38286 21128 38292 21140
rect 38247 21100 38292 21128
rect 36817 21091 36875 21097
rect 38286 21088 38292 21100
rect 38344 21088 38350 21140
rect 35713 21063 35771 21069
rect 35713 21060 35725 21063
rect 25056 21032 35725 21060
rect 35713 21029 35725 21032
rect 35759 21029 35771 21063
rect 35713 21023 35771 21029
rect 35802 21020 35808 21072
rect 35860 21060 35866 21072
rect 35860 21032 36860 21060
rect 35860 21020 35866 21032
rect 19518 20992 19524 21004
rect 18708 20964 19380 20992
rect 19479 20964 19524 20992
rect 18708 20936 18736 20964
rect 19518 20952 19524 20964
rect 19576 20952 19582 21004
rect 28074 20992 28080 21004
rect 25424 20964 28080 20992
rect 1940 20927 1998 20933
rect 1940 20893 1952 20927
rect 1986 20924 1998 20927
rect 2222 20924 2228 20936
rect 1986 20896 2228 20924
rect 1986 20893 1998 20896
rect 1940 20887 1998 20893
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 7006 20884 7012 20936
rect 7064 20924 7070 20936
rect 7653 20927 7711 20933
rect 7653 20924 7665 20927
rect 7064 20896 7665 20924
rect 7064 20884 7070 20896
rect 7653 20893 7665 20896
rect 7699 20924 7711 20927
rect 7742 20924 7748 20936
rect 7699 20896 7748 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 7742 20884 7748 20896
rect 7800 20884 7806 20936
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 8021 20927 8079 20933
rect 7892 20896 7985 20924
rect 8021 20912 8033 20927
rect 8067 20912 8079 20927
rect 10502 20924 10508 20936
rect 7892 20884 7898 20896
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 7852 20856 7880 20884
rect 8018 20860 8024 20912
rect 8076 20860 8082 20912
rect 10463 20896 10508 20924
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 15838 20924 15844 20936
rect 15751 20896 15844 20924
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 17494 20924 17500 20936
rect 17455 20896 17500 20924
rect 16117 20887 16175 20893
rect 7616 20828 7880 20856
rect 7616 20816 7622 20828
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 13173 20859 13231 20865
rect 13173 20856 13185 20859
rect 12492 20828 13185 20856
rect 12492 20816 12498 20828
rect 13173 20825 13185 20828
rect 13219 20856 13231 20859
rect 13722 20856 13728 20868
rect 13219 20828 13728 20856
rect 13219 20825 13231 20828
rect 13173 20819 13231 20825
rect 13722 20816 13728 20828
rect 13780 20816 13786 20868
rect 2958 20748 2964 20800
rect 3016 20788 3022 20800
rect 3053 20791 3111 20797
rect 3053 20788 3065 20791
rect 3016 20760 3065 20788
rect 3016 20748 3022 20760
rect 3053 20757 3065 20760
rect 3099 20788 3111 20791
rect 6914 20788 6920 20800
rect 3099 20760 6920 20788
rect 3099 20757 3111 20760
rect 3053 20751 3111 20757
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 7285 20791 7343 20797
rect 7285 20757 7297 20791
rect 7331 20788 7343 20791
rect 8662 20788 8668 20800
rect 7331 20760 8668 20788
rect 7331 20757 7343 20760
rect 7285 20751 7343 20757
rect 8662 20748 8668 20760
rect 8720 20748 8726 20800
rect 10321 20791 10379 20797
rect 10321 20757 10333 20791
rect 10367 20788 10379 20791
rect 10686 20788 10692 20800
rect 10367 20760 10692 20788
rect 10367 20757 10379 20760
rect 10321 20751 10379 20757
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 11112 20760 13277 20788
rect 11112 20748 11118 20760
rect 13265 20757 13277 20760
rect 13311 20788 13323 20791
rect 15562 20788 15568 20800
rect 13311 20760 15568 20788
rect 13311 20757 13323 20760
rect 13265 20751 13323 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 15856 20788 15884 20884
rect 16132 20856 16160 20887
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 17678 20924 17684 20936
rect 17639 20896 17684 20924
rect 17678 20884 17684 20896
rect 17736 20924 17742 20936
rect 18690 20924 18696 20936
rect 17736 20896 18696 20924
rect 17736 20884 17742 20896
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 19288 20884 19294 20936
rect 19346 20924 19352 20936
rect 19403 20927 19461 20933
rect 19403 20924 19415 20927
rect 19346 20896 19415 20924
rect 19346 20884 19352 20896
rect 19403 20893 19415 20896
rect 19449 20893 19461 20927
rect 19614 20927 19672 20933
rect 19614 20900 19626 20927
rect 19403 20887 19461 20893
rect 19505 20893 19626 20900
rect 19660 20893 19672 20927
rect 19505 20887 19672 20893
rect 19505 20872 19657 20887
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 21545 20927 21603 20933
rect 19760 20896 19805 20924
rect 19760 20884 19766 20896
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 21634 20924 21640 20936
rect 21591 20896 21640 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 21634 20884 21640 20896
rect 21692 20884 21698 20936
rect 25424 20933 25452 20964
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 28258 20952 28264 21004
rect 28316 20992 28322 21004
rect 32582 20992 32588 21004
rect 28316 20964 32444 20992
rect 32543 20964 32588 20992
rect 28316 20952 28322 20964
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20924 25743 20927
rect 25774 20924 25780 20936
rect 25731 20896 25780 20924
rect 25731 20893 25743 20896
rect 25685 20887 25743 20893
rect 25774 20884 25780 20896
rect 25832 20924 25838 20936
rect 26234 20924 26240 20936
rect 25832 20896 26240 20924
rect 25832 20884 25838 20896
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26712 20896 27384 20924
rect 18138 20856 18144 20868
rect 16132 20828 18144 20856
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 19208 20828 19334 20856
rect 19208 20816 19214 20828
rect 17862 20788 17868 20800
rect 15856 20760 17868 20788
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 19306 20788 19334 20828
rect 19505 20788 19533 20872
rect 21812 20859 21870 20865
rect 21812 20825 21824 20859
rect 21858 20856 21870 20859
rect 22002 20856 22008 20868
rect 21858 20828 22008 20856
rect 21858 20825 21870 20828
rect 21812 20819 21870 20825
rect 22002 20816 22008 20828
rect 22060 20816 22066 20868
rect 23014 20816 23020 20868
rect 23072 20856 23078 20868
rect 26712 20856 26740 20896
rect 23072 20828 26740 20856
rect 23072 20816 23078 20828
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 27246 20856 27252 20868
rect 26844 20828 27252 20856
rect 26844 20816 26850 20828
rect 27246 20816 27252 20828
rect 27304 20816 27310 20868
rect 27356 20856 27384 20896
rect 27614 20884 27620 20936
rect 27672 20924 27678 20936
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 27672 20896 28181 20924
rect 27672 20884 27678 20896
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 28169 20887 28227 20893
rect 31570 20884 31576 20936
rect 31628 20924 31634 20936
rect 32309 20927 32367 20933
rect 32309 20924 32321 20927
rect 31628 20896 32321 20924
rect 31628 20884 31634 20896
rect 32309 20893 32321 20896
rect 32355 20893 32367 20927
rect 32416 20924 32444 20964
rect 32582 20952 32588 20964
rect 32640 20952 32646 21004
rect 32766 20952 32772 21004
rect 32824 20992 32830 21004
rect 32824 20964 35204 20992
rect 32824 20952 32830 20964
rect 33594 20924 33600 20936
rect 32416 20896 33600 20924
rect 32309 20887 32367 20893
rect 33594 20884 33600 20896
rect 33652 20884 33658 20936
rect 34698 20884 34704 20936
rect 34756 20924 34762 20936
rect 35176 20933 35204 20964
rect 35069 20927 35127 20933
rect 35069 20924 35081 20927
rect 34756 20896 35081 20924
rect 34756 20884 34762 20896
rect 35069 20893 35081 20896
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35162 20927 35220 20933
rect 35162 20893 35174 20927
rect 35208 20893 35220 20927
rect 35162 20887 35220 20893
rect 35534 20927 35592 20933
rect 35534 20893 35546 20927
rect 35580 20924 35592 20927
rect 35580 20896 35664 20924
rect 35580 20893 35592 20896
rect 35534 20887 35592 20893
rect 34238 20856 34244 20868
rect 27356 20828 34244 20856
rect 34238 20816 34244 20828
rect 34296 20816 34302 20868
rect 19306 20760 19533 20788
rect 22370 20748 22376 20800
rect 22428 20788 22434 20800
rect 22925 20791 22983 20797
rect 22925 20788 22937 20791
rect 22428 20760 22937 20788
rect 22428 20748 22434 20760
rect 22925 20757 22937 20760
rect 22971 20757 22983 20791
rect 22925 20751 22983 20757
rect 23382 20748 23388 20800
rect 23440 20788 23446 20800
rect 25593 20791 25651 20797
rect 25593 20788 25605 20791
rect 23440 20760 25605 20788
rect 23440 20748 23446 20760
rect 25593 20757 25605 20760
rect 25639 20788 25651 20791
rect 26050 20788 26056 20800
rect 25639 20760 26056 20788
rect 25639 20757 25651 20760
rect 25593 20751 25651 20757
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 27341 20791 27399 20797
rect 27341 20757 27353 20791
rect 27387 20788 27399 20791
rect 27522 20788 27528 20800
rect 27387 20760 27528 20788
rect 27387 20757 27399 20760
rect 27341 20751 27399 20757
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 27982 20788 27988 20800
rect 27943 20760 27988 20788
rect 27982 20748 27988 20760
rect 28040 20748 28046 20800
rect 28074 20748 28080 20800
rect 28132 20788 28138 20800
rect 34790 20788 34796 20800
rect 28132 20760 34796 20788
rect 28132 20748 28138 20760
rect 34790 20748 34796 20760
rect 34848 20748 34854 20800
rect 35091 20788 35119 20887
rect 35342 20856 35348 20868
rect 35303 20828 35348 20856
rect 35342 20816 35348 20828
rect 35400 20816 35406 20868
rect 35434 20816 35440 20868
rect 35492 20856 35498 20868
rect 35636 20856 35664 20896
rect 35802 20884 35808 20936
rect 35860 20924 35866 20936
rect 36173 20927 36231 20933
rect 36173 20924 36185 20927
rect 35860 20896 36185 20924
rect 35860 20884 35866 20896
rect 36173 20893 36185 20896
rect 36219 20893 36231 20927
rect 36173 20887 36231 20893
rect 36262 20884 36268 20936
rect 36320 20924 36326 20936
rect 36638 20927 36696 20933
rect 36320 20896 36365 20924
rect 36320 20884 36326 20896
rect 36638 20893 36650 20927
rect 36684 20924 36696 20927
rect 36832 20924 36860 21032
rect 38473 20927 38531 20933
rect 38473 20924 38485 20927
rect 36684 20896 36768 20924
rect 36832 20896 38485 20924
rect 36684 20893 36696 20896
rect 36638 20887 36696 20893
rect 35492 20828 35537 20856
rect 35636 20828 36216 20856
rect 35492 20816 35498 20828
rect 36188 20800 36216 20828
rect 36354 20816 36360 20868
rect 36412 20856 36418 20868
rect 36449 20859 36507 20865
rect 36449 20856 36461 20859
rect 36412 20828 36461 20856
rect 36412 20816 36418 20828
rect 36449 20825 36461 20828
rect 36495 20825 36507 20859
rect 36449 20819 36507 20825
rect 36538 20816 36544 20868
rect 36596 20856 36602 20868
rect 36596 20828 36641 20856
rect 36596 20816 36602 20828
rect 35802 20788 35808 20800
rect 35091 20760 35808 20788
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 36170 20748 36176 20800
rect 36228 20788 36234 20800
rect 36740 20788 36768 20896
rect 38473 20893 38485 20896
rect 38519 20893 38531 20927
rect 38746 20924 38752 20936
rect 38707 20896 38752 20924
rect 38473 20887 38531 20893
rect 38746 20884 38752 20896
rect 38804 20884 38810 20936
rect 37826 20816 37832 20868
rect 37884 20856 37890 20868
rect 38657 20859 38715 20865
rect 38657 20856 38669 20859
rect 37884 20828 38669 20856
rect 37884 20816 37890 20828
rect 38657 20825 38669 20828
rect 38703 20856 38715 20859
rect 39850 20856 39856 20868
rect 38703 20828 39856 20856
rect 38703 20825 38715 20828
rect 38657 20819 38715 20825
rect 39850 20816 39856 20828
rect 39908 20816 39914 20868
rect 36228 20760 36768 20788
rect 36228 20748 36234 20760
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 2133 20587 2191 20593
rect 2133 20553 2145 20587
rect 2179 20584 2191 20587
rect 2406 20584 2412 20596
rect 2179 20556 2412 20584
rect 2179 20553 2191 20556
rect 2133 20547 2191 20553
rect 2406 20544 2412 20556
rect 2464 20544 2470 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 2958 20584 2964 20596
rect 2547 20556 2964 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 7193 20587 7251 20593
rect 7193 20553 7205 20587
rect 7239 20584 7251 20587
rect 8018 20584 8024 20596
rect 7239 20556 8024 20584
rect 7239 20553 7251 20556
rect 7193 20547 7251 20553
rect 8018 20544 8024 20556
rect 8076 20544 8082 20596
rect 10229 20587 10287 20593
rect 10229 20553 10241 20587
rect 10275 20584 10287 20587
rect 10502 20584 10508 20596
rect 10275 20556 10508 20584
rect 10275 20553 10287 20556
rect 10229 20547 10287 20553
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10597 20587 10655 20593
rect 10597 20553 10609 20587
rect 10643 20584 10655 20587
rect 11054 20584 11060 20596
rect 10643 20556 11060 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 17957 20587 18015 20593
rect 17957 20553 17969 20587
rect 18003 20584 18015 20587
rect 19288 20584 19294 20596
rect 18003 20556 19294 20584
rect 18003 20553 18015 20556
rect 17957 20547 18015 20553
rect 19288 20544 19294 20556
rect 19346 20544 19352 20596
rect 19720 20556 20116 20584
rect 8110 20516 8116 20528
rect 7024 20488 8116 20516
rect 7024 20460 7052 20488
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 12894 20516 12900 20528
rect 12492 20488 12537 20516
rect 12855 20488 12900 20516
rect 12492 20476 12498 20488
rect 12894 20476 12900 20488
rect 12952 20476 12958 20528
rect 13081 20519 13139 20525
rect 13081 20485 13093 20519
rect 13127 20516 13139 20519
rect 13170 20516 13176 20528
rect 13127 20488 13176 20516
rect 13127 20485 13139 20488
rect 13081 20479 13139 20485
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 16942 20476 16948 20528
rect 17000 20516 17006 20528
rect 19720 20516 19748 20556
rect 17000 20488 19748 20516
rect 20088 20516 20116 20556
rect 20162 20544 20168 20596
rect 20220 20584 20226 20596
rect 22370 20584 22376 20596
rect 20220 20556 22232 20584
rect 22331 20556 22376 20584
rect 20220 20544 20226 20556
rect 21726 20516 21732 20528
rect 20088 20488 21732 20516
rect 17000 20476 17006 20488
rect 21726 20476 21732 20488
rect 21784 20476 21790 20528
rect 22002 20516 22008 20528
rect 21963 20488 22008 20516
rect 22002 20476 22008 20488
rect 22060 20476 22066 20528
rect 22204 20516 22232 20556
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 25774 20584 25780 20596
rect 25735 20556 25780 20584
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 27525 20587 27583 20593
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 27614 20584 27620 20596
rect 27571 20556 27620 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 27614 20544 27620 20556
rect 27672 20544 27678 20596
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 34054 20584 34060 20596
rect 27764 20556 34060 20584
rect 27764 20544 27770 20556
rect 34054 20544 34060 20556
rect 34112 20544 34118 20596
rect 36354 20584 36360 20596
rect 36004 20556 36360 20584
rect 22204 20488 27844 20516
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20417 1455 20451
rect 1397 20411 1455 20417
rect 1412 20312 1440 20411
rect 3326 20408 3332 20460
rect 3384 20448 3390 20460
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3384 20420 3801 20448
rect 3384 20408 3390 20420
rect 3789 20417 3801 20420
rect 3835 20417 3847 20451
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 3789 20411 3847 20417
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7006 20448 7012 20460
rect 6967 20420 7012 20448
rect 7006 20408 7012 20420
rect 7064 20408 7070 20460
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20448 7711 20451
rect 7834 20448 7840 20460
rect 7699 20420 7840 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 8846 20448 8852 20460
rect 7975 20420 8852 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 8846 20408 8852 20420
rect 8904 20408 8910 20460
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12253 20451 12311 20457
rect 12253 20448 12265 20451
rect 11848 20420 12265 20448
rect 11848 20408 11854 20420
rect 12253 20417 12265 20420
rect 12299 20417 12311 20451
rect 12253 20411 12311 20417
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 16574 20448 16580 20460
rect 15611 20420 16580 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 16574 20408 16580 20420
rect 16632 20408 16638 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17126 20448 17132 20460
rect 16715 20420 17132 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 18046 20448 18052 20460
rect 17604 20420 18052 20448
rect 2590 20380 2596 20392
rect 2551 20352 2596 20380
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 2682 20340 2688 20392
rect 2740 20380 2746 20392
rect 7742 20380 7748 20392
rect 2740 20352 2785 20380
rect 7703 20352 7748 20380
rect 2740 20340 2746 20352
rect 7742 20340 7748 20352
rect 7800 20340 7806 20392
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10468 20352 10701 20380
rect 10468 20340 10474 20352
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20380 15347 20383
rect 15470 20380 15476 20392
rect 15335 20352 15476 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 9674 20312 9680 20324
rect 1412 20284 9680 20312
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 10594 20312 10600 20324
rect 9916 20284 10600 20312
rect 9916 20272 9922 20284
rect 10594 20272 10600 20284
rect 10652 20312 10658 20324
rect 10796 20312 10824 20343
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16945 20383 17003 20389
rect 16945 20349 16957 20383
rect 16991 20380 17003 20383
rect 17604 20380 17632 20420
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 19242 20408 19248 20460
rect 19300 20448 19306 20460
rect 19334 20448 19340 20460
rect 19300 20410 19340 20448
rect 19300 20408 19306 20410
rect 19334 20408 19340 20410
rect 19392 20408 19398 20460
rect 19812 20457 20024 20470
rect 19797 20451 20024 20457
rect 19797 20417 19809 20451
rect 19843 20448 20024 20451
rect 19843 20442 22140 20448
rect 19843 20417 19855 20442
rect 19996 20420 22140 20442
rect 19797 20411 19855 20417
rect 16991 20352 17632 20380
rect 16991 20349 17003 20352
rect 16945 20343 17003 20349
rect 17862 20340 17868 20392
rect 17920 20380 17926 20392
rect 18141 20383 18199 20389
rect 18141 20380 18153 20383
rect 17920 20352 18153 20380
rect 17920 20340 17926 20352
rect 18141 20349 18153 20352
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 18233 20383 18291 20389
rect 18233 20349 18245 20383
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20349 18383 20383
rect 18325 20343 18383 20349
rect 10652 20284 10824 20312
rect 10652 20272 10658 20284
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15102 20312 15108 20324
rect 14884 20284 15108 20312
rect 14884 20272 14890 20284
rect 15102 20272 15108 20284
rect 15160 20272 15166 20324
rect 15562 20272 15568 20324
rect 15620 20312 15626 20324
rect 17954 20312 17960 20324
rect 15620 20284 17960 20312
rect 15620 20272 15626 20284
rect 17954 20272 17960 20284
rect 18012 20312 18018 20324
rect 18248 20312 18276 20343
rect 18012 20284 18276 20312
rect 18340 20312 18368 20343
rect 18414 20340 18420 20392
rect 18472 20380 18478 20392
rect 19518 20380 19524 20392
rect 18472 20352 18517 20380
rect 19479 20352 19524 20380
rect 18472 20340 18478 20352
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 19886 20380 19892 20392
rect 19760 20352 19805 20380
rect 19847 20352 19892 20380
rect 19760 20340 19766 20352
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20070 20380 20076 20392
rect 20027 20352 20076 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20070 20340 20076 20352
rect 20128 20340 20134 20392
rect 22112 20380 22140 20420
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22462 20448 22468 20460
rect 22244 20420 22289 20448
rect 22423 20420 22468 20448
rect 22244 20408 22250 20420
rect 22462 20408 22468 20420
rect 22520 20408 22526 20460
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20448 25743 20451
rect 26142 20448 26148 20460
rect 25731 20420 26148 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 27154 20448 27160 20460
rect 27115 20420 27160 20448
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 27338 20448 27344 20460
rect 27299 20420 27344 20448
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27816 20448 27844 20488
rect 27982 20476 27988 20528
rect 28040 20516 28046 20528
rect 28230 20519 28288 20525
rect 28230 20516 28242 20519
rect 28040 20488 28242 20516
rect 28040 20476 28046 20488
rect 28230 20485 28242 20488
rect 28276 20485 28288 20519
rect 28230 20479 28288 20485
rect 35342 20476 35348 20528
rect 35400 20516 35406 20528
rect 36004 20525 36032 20556
rect 36354 20544 36360 20556
rect 36412 20544 36418 20596
rect 35989 20519 36047 20525
rect 35989 20516 36001 20519
rect 35400 20488 36001 20516
rect 35400 20476 35406 20488
rect 35989 20485 36001 20488
rect 36035 20485 36047 20519
rect 35989 20479 36047 20485
rect 36081 20519 36139 20525
rect 36081 20485 36093 20519
rect 36127 20516 36139 20519
rect 36446 20516 36452 20528
rect 36127 20488 36452 20516
rect 36127 20485 36139 20488
rect 36081 20479 36139 20485
rect 36446 20476 36452 20488
rect 36504 20476 36510 20528
rect 34790 20448 34796 20460
rect 27816 20420 34796 20448
rect 34790 20408 34796 20420
rect 34848 20408 34854 20460
rect 35710 20448 35716 20460
rect 35671 20420 35716 20448
rect 35710 20408 35716 20420
rect 35768 20408 35774 20460
rect 35861 20451 35919 20457
rect 35861 20417 35873 20451
rect 35907 20448 35919 20451
rect 35907 20420 36124 20448
rect 35907 20417 35919 20420
rect 35861 20411 35919 20417
rect 27706 20380 27712 20392
rect 22112 20352 27712 20380
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 27890 20340 27896 20392
rect 27948 20380 27954 20392
rect 27985 20383 28043 20389
rect 27985 20380 27997 20383
rect 27948 20352 27997 20380
rect 27948 20340 27954 20352
rect 27985 20349 27997 20352
rect 28031 20349 28043 20383
rect 36096 20380 36124 20420
rect 36170 20408 36176 20460
rect 36228 20457 36234 20460
rect 36228 20448 36236 20457
rect 36228 20420 36273 20448
rect 36228 20411 36236 20420
rect 36228 20408 36234 20411
rect 38746 20408 38752 20460
rect 38804 20448 38810 20460
rect 39373 20451 39431 20457
rect 39373 20448 39385 20451
rect 38804 20420 39385 20448
rect 38804 20408 38810 20420
rect 39373 20417 39385 20420
rect 39419 20417 39431 20451
rect 39373 20411 39431 20417
rect 38194 20380 38200 20392
rect 36096 20352 38200 20380
rect 27985 20343 28043 20349
rect 38194 20340 38200 20352
rect 38252 20340 38258 20392
rect 39114 20380 39120 20392
rect 39075 20352 39120 20380
rect 39114 20340 39120 20352
rect 39172 20340 39178 20392
rect 23382 20312 23388 20324
rect 18340 20284 23388 20312
rect 18012 20272 18018 20284
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 36357 20315 36415 20321
rect 36357 20312 36369 20315
rect 28966 20284 36369 20312
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 3602 20244 3608 20256
rect 3563 20216 3608 20244
rect 3602 20204 3608 20216
rect 3660 20204 3666 20256
rect 7650 20244 7656 20256
rect 7611 20216 7656 20244
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 9582 20244 9588 20256
rect 8159 20216 9588 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 13078 20244 13084 20256
rect 13039 20216 13084 20244
rect 13078 20204 13084 20216
rect 13136 20204 13142 20256
rect 13265 20247 13323 20253
rect 13265 20213 13277 20247
rect 13311 20244 13323 20247
rect 20346 20244 20352 20256
rect 13311 20216 20352 20244
rect 13311 20213 13323 20216
rect 13265 20207 13323 20213
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 28966 20244 28994 20284
rect 36357 20281 36369 20284
rect 36403 20281 36415 20315
rect 36357 20275 36415 20281
rect 21784 20216 28994 20244
rect 29365 20247 29423 20253
rect 21784 20204 21790 20216
rect 29365 20213 29377 20247
rect 29411 20244 29423 20247
rect 29546 20244 29552 20256
rect 29411 20216 29552 20244
rect 29411 20213 29423 20216
rect 29365 20207 29423 20213
rect 29546 20204 29552 20216
rect 29604 20204 29610 20256
rect 40034 20204 40040 20256
rect 40092 20244 40098 20256
rect 40497 20247 40555 20253
rect 40497 20244 40509 20247
rect 40092 20216 40509 20244
rect 40092 20204 40098 20216
rect 40497 20213 40509 20216
rect 40543 20213 40555 20247
rect 40497 20207 40555 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 2501 20043 2559 20049
rect 2501 20009 2513 20043
rect 2547 20040 2559 20043
rect 2590 20040 2596 20052
rect 2547 20012 2596 20040
rect 2547 20009 2559 20012
rect 2501 20003 2559 20009
rect 2590 20000 2596 20012
rect 2648 20000 2654 20052
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 7377 20043 7435 20049
rect 3476 20012 4752 20040
rect 3476 20000 3482 20012
rect 4724 19972 4752 20012
rect 7377 20009 7389 20043
rect 7423 20040 7435 20043
rect 8294 20040 8300 20052
rect 7423 20012 8300 20040
rect 7423 20009 7435 20012
rect 7377 20003 7435 20009
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 11790 20040 11796 20052
rect 11751 20012 11796 20040
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 12894 20040 12900 20052
rect 12851 20012 12900 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 14645 20043 14703 20049
rect 14645 20009 14657 20043
rect 14691 20040 14703 20043
rect 15930 20040 15936 20052
rect 14691 20012 15936 20040
rect 14691 20009 14703 20012
rect 14645 20003 14703 20009
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 24118 20040 24124 20052
rect 17552 20012 24124 20040
rect 17552 20000 17558 20012
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 27154 20000 27160 20052
rect 27212 20040 27218 20052
rect 28629 20043 28687 20049
rect 28629 20040 28641 20043
rect 27212 20012 28641 20040
rect 27212 20000 27218 20012
rect 28629 20009 28641 20012
rect 28675 20009 28687 20043
rect 38746 20040 38752 20052
rect 28629 20003 28687 20009
rect 28736 20012 38424 20040
rect 38707 20012 38752 20040
rect 23014 19972 23020 19984
rect 4724 19944 8524 19972
rect 1486 19864 1492 19916
rect 1544 19904 1550 19916
rect 3789 19907 3847 19913
rect 3789 19904 3801 19907
rect 1544 19876 3801 19904
rect 1544 19864 1550 19876
rect 3789 19873 3801 19876
rect 3835 19873 3847 19907
rect 3789 19867 3847 19873
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 7285 19907 7343 19913
rect 7285 19904 7297 19907
rect 6880 19876 7297 19904
rect 6880 19864 6886 19876
rect 7285 19873 7297 19876
rect 7331 19904 7343 19907
rect 8389 19907 8447 19913
rect 8389 19904 8401 19907
rect 7331 19876 8401 19904
rect 7331 19873 7343 19876
rect 7285 19867 7343 19873
rect 8389 19873 8401 19876
rect 8435 19873 8447 19907
rect 8389 19867 8447 19873
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 2774 19836 2780 19848
rect 2731 19808 2780 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 3602 19796 3608 19848
rect 3660 19836 3666 19848
rect 4045 19839 4103 19845
rect 4045 19836 4057 19839
rect 3660 19808 4057 19836
rect 3660 19796 3666 19808
rect 4045 19805 4057 19808
rect 4091 19805 4103 19839
rect 4045 19799 4103 19805
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7156 19808 7389 19836
rect 7156 19796 7162 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 7926 19836 7932 19848
rect 7377 19799 7435 19805
rect 7484 19808 7932 19836
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 2041 19771 2099 19777
rect 2041 19737 2053 19771
rect 2087 19768 2099 19771
rect 2130 19768 2136 19780
rect 2087 19740 2136 19768
rect 2087 19737 2099 19740
rect 2041 19731 2099 19737
rect 2130 19728 2136 19740
rect 2188 19728 2194 19780
rect 6914 19768 6920 19780
rect 6827 19740 6920 19768
rect 6914 19728 6920 19740
rect 6972 19768 6978 19780
rect 7484 19768 7512 19808
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 8018 19768 8024 19780
rect 6972 19740 7512 19768
rect 7979 19740 8024 19768
rect 6972 19728 6978 19740
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 8110 19728 8116 19780
rect 8168 19768 8174 19780
rect 8205 19771 8263 19777
rect 8205 19768 8217 19771
rect 8168 19740 8217 19768
rect 8168 19728 8174 19740
rect 8205 19737 8217 19740
rect 8251 19737 8263 19771
rect 8496 19768 8524 19944
rect 13556 19944 15705 19972
rect 10226 19864 10232 19916
rect 10284 19904 10290 19916
rect 13556 19913 13584 19944
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 10284 19876 10425 19904
rect 10284 19864 10290 19876
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19873 13599 19907
rect 13541 19867 13599 19873
rect 13722 19864 13728 19916
rect 13780 19904 13786 19916
rect 15562 19904 15568 19916
rect 13780 19876 15568 19904
rect 13780 19864 13786 19876
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 15677 19904 15705 19944
rect 16408 19944 23020 19972
rect 16408 19904 16436 19944
rect 23014 19932 23020 19944
rect 23072 19932 23078 19984
rect 18414 19904 18420 19916
rect 15677 19876 16436 19904
rect 16776 19876 18420 19904
rect 10686 19845 10692 19848
rect 10680 19836 10692 19845
rect 10647 19808 10692 19836
rect 10680 19799 10692 19808
rect 10686 19796 10692 19799
rect 10744 19796 10750 19848
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 13078 19796 13084 19808
rect 13136 19836 13142 19848
rect 13630 19836 13636 19848
rect 13136 19808 13636 19836
rect 13136 19796 13142 19808
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 15378 19836 15384 19848
rect 14660 19808 15384 19836
rect 14660 19777 14688 19808
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19836 15807 19839
rect 15930 19836 15936 19848
rect 15795 19808 15936 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 12989 19771 13047 19777
rect 12989 19768 13001 19771
rect 8496 19740 13001 19768
rect 8205 19731 8263 19737
rect 12989 19737 13001 19740
rect 13035 19737 13047 19771
rect 12989 19731 13047 19737
rect 14461 19771 14519 19777
rect 14461 19737 14473 19771
rect 14507 19737 14519 19771
rect 14660 19771 14719 19777
rect 14660 19740 14673 19771
rect 14461 19731 14519 19737
rect 14661 19737 14673 19740
rect 14707 19737 14719 19771
rect 14661 19731 14719 19737
rect 14752 19740 15424 19768
rect 5166 19700 5172 19712
rect 5127 19672 5172 19700
rect 5166 19660 5172 19672
rect 5224 19700 5230 19712
rect 7006 19700 7012 19712
rect 5224 19672 7012 19700
rect 5224 19660 5230 19672
rect 7006 19660 7012 19672
rect 7064 19660 7070 19712
rect 7561 19703 7619 19709
rect 7561 19669 7573 19703
rect 7607 19700 7619 19703
rect 7926 19700 7932 19712
rect 7607 19672 7932 19700
rect 7607 19669 7619 19672
rect 7561 19663 7619 19669
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 14476 19700 14504 19731
rect 14752 19700 14780 19740
rect 15396 19712 15424 19740
rect 14476 19672 14780 19700
rect 14829 19703 14887 19709
rect 14829 19669 14841 19703
rect 14875 19700 14887 19703
rect 15102 19700 15108 19712
rect 14875 19672 15108 19700
rect 14875 19669 14887 19672
rect 14829 19663 14887 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15378 19660 15384 19712
rect 15436 19660 15442 19712
rect 15488 19700 15516 19799
rect 15562 19728 15568 19780
rect 15620 19768 15626 19780
rect 15672 19768 15700 19799
rect 15930 19796 15936 19808
rect 15988 19836 15994 19848
rect 16776 19836 16804 19876
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 19702 19904 19708 19916
rect 19663 19876 19708 19904
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 19794 19864 19800 19916
rect 19852 19904 19858 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19852 19876 19993 19904
rect 19852 19864 19858 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20165 19907 20223 19913
rect 20165 19873 20177 19907
rect 20211 19904 20223 19907
rect 20254 19904 20260 19916
rect 20211 19876 20260 19904
rect 20211 19873 20223 19876
rect 20165 19867 20223 19873
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 22186 19864 22192 19916
rect 22244 19904 22250 19916
rect 22462 19904 22468 19916
rect 22244 19876 22468 19904
rect 22244 19864 22250 19876
rect 22462 19864 22468 19876
rect 22520 19904 22526 19916
rect 28736 19904 28764 20012
rect 28902 19932 28908 19984
rect 28960 19972 28966 19984
rect 38289 19975 38347 19981
rect 28960 19944 30880 19972
rect 28960 19932 28966 19944
rect 22520 19876 24532 19904
rect 22520 19864 22526 19876
rect 17402 19836 17408 19848
rect 15988 19808 16804 19836
rect 17363 19808 17408 19836
rect 15988 19796 15994 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 19886 19836 19892 19848
rect 19847 19808 19892 19836
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19836 20131 19839
rect 20119 19808 20300 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 15620 19740 15700 19768
rect 15620 19728 15626 19740
rect 16114 19728 16120 19780
rect 16172 19768 16178 19780
rect 20162 19768 20168 19780
rect 16172 19740 20168 19768
rect 16172 19728 16178 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 15838 19700 15844 19712
rect 15488 19672 15844 19700
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 20272 19700 20300 19808
rect 21634 19796 21640 19848
rect 21692 19836 21698 19848
rect 24394 19836 24400 19848
rect 21692 19808 24400 19836
rect 21692 19796 21698 19808
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 24504 19836 24532 19876
rect 25424 19876 28764 19904
rect 25424 19836 25452 19876
rect 28994 19864 29000 19916
rect 29052 19904 29058 19916
rect 29641 19907 29699 19913
rect 29641 19904 29653 19907
rect 29052 19876 29653 19904
rect 29052 19864 29058 19876
rect 29641 19873 29653 19876
rect 29687 19873 29699 19907
rect 29641 19867 29699 19873
rect 29730 19864 29736 19916
rect 29788 19904 29794 19916
rect 29825 19907 29883 19913
rect 29825 19904 29837 19907
rect 29788 19876 29837 19904
rect 29788 19864 29794 19876
rect 29825 19873 29837 19876
rect 29871 19873 29883 19907
rect 29825 19867 29883 19873
rect 24504 19808 25452 19836
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19805 28687 19839
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 28629 19799 28687 19805
rect 20346 19728 20352 19780
rect 20404 19768 20410 19780
rect 22370 19768 22376 19780
rect 20404 19740 22376 19768
rect 20404 19728 20410 19740
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 24670 19777 24676 19780
rect 24664 19731 24676 19777
rect 24728 19768 24734 19780
rect 24728 19740 24764 19768
rect 24670 19728 24676 19731
rect 24728 19728 24734 19740
rect 26234 19728 26240 19780
rect 26292 19768 26298 19780
rect 27154 19768 27160 19780
rect 26292 19740 27160 19768
rect 26292 19728 26298 19740
rect 27154 19728 27160 19740
rect 27212 19728 27218 19780
rect 27249 19771 27307 19777
rect 27249 19737 27261 19771
rect 27295 19768 27307 19771
rect 27522 19768 27528 19780
rect 27295 19740 27528 19768
rect 27295 19737 27307 19740
rect 27249 19731 27307 19737
rect 27522 19728 27528 19740
rect 27580 19728 27586 19780
rect 28644 19768 28672 19799
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 29546 19836 29552 19848
rect 29507 19808 29552 19836
rect 29546 19796 29552 19808
rect 29604 19836 29610 19848
rect 30558 19836 30564 19848
rect 29604 19808 30564 19836
rect 29604 19796 29610 19808
rect 30558 19796 30564 19808
rect 30616 19796 30622 19848
rect 30742 19836 30748 19848
rect 30703 19808 30748 19836
rect 30742 19796 30748 19808
rect 30800 19796 30806 19848
rect 30852 19836 30880 19944
rect 38289 19941 38301 19975
rect 38335 19941 38347 19975
rect 38396 19972 38424 20012
rect 38746 20000 38752 20012
rect 38804 20000 38810 20052
rect 39114 20000 39120 20052
rect 39172 20040 39178 20052
rect 40494 20040 40500 20052
rect 39172 20012 40500 20040
rect 39172 20000 39178 20012
rect 40494 20000 40500 20012
rect 40552 20000 40558 20052
rect 38396 19944 39252 19972
rect 38289 19935 38347 19941
rect 31202 19904 31208 19916
rect 31163 19876 31208 19904
rect 31202 19864 31208 19876
rect 31260 19864 31266 19916
rect 38304 19904 38332 19935
rect 38838 19904 38844 19916
rect 36188 19876 38240 19904
rect 38304 19876 38844 19904
rect 35802 19836 35808 19848
rect 30852 19808 34192 19836
rect 35763 19808 35808 19836
rect 29825 19771 29883 19777
rect 29825 19768 29837 19771
rect 28644 19740 29837 19768
rect 29825 19737 29837 19740
rect 29871 19737 29883 19771
rect 31450 19771 31508 19777
rect 31450 19768 31462 19771
rect 29825 19731 29883 19737
rect 30760 19740 31462 19768
rect 25038 19700 25044 19712
rect 20272 19672 25044 19700
rect 25038 19660 25044 19672
rect 25096 19700 25102 19712
rect 25777 19703 25835 19709
rect 25777 19700 25789 19703
rect 25096 19672 25789 19700
rect 25096 19660 25102 19672
rect 25777 19669 25789 19672
rect 25823 19669 25835 19703
rect 25777 19663 25835 19669
rect 26142 19660 26148 19712
rect 26200 19700 26206 19712
rect 27341 19703 27399 19709
rect 27341 19700 27353 19703
rect 26200 19672 27353 19700
rect 26200 19660 26206 19672
rect 27341 19669 27353 19672
rect 27387 19669 27399 19703
rect 27540 19700 27568 19728
rect 29086 19700 29092 19712
rect 27540 19672 29092 19700
rect 27341 19663 27399 19669
rect 29086 19660 29092 19672
rect 29144 19700 29150 19712
rect 29730 19700 29736 19712
rect 29144 19672 29736 19700
rect 29144 19660 29150 19672
rect 29730 19660 29736 19672
rect 29788 19700 29794 19712
rect 30098 19700 30104 19712
rect 29788 19672 30104 19700
rect 29788 19660 29794 19672
rect 30098 19660 30104 19672
rect 30156 19660 30162 19712
rect 30561 19703 30619 19709
rect 30561 19669 30573 19703
rect 30607 19700 30619 19703
rect 30760 19700 30788 19740
rect 31450 19737 31462 19740
rect 31496 19737 31508 19771
rect 31450 19731 31508 19737
rect 32582 19700 32588 19712
rect 30607 19672 30788 19700
rect 32543 19672 32588 19700
rect 30607 19669 30619 19672
rect 30561 19663 30619 19669
rect 32582 19660 32588 19672
rect 32640 19660 32646 19712
rect 34164 19700 34192 19808
rect 35802 19796 35808 19808
rect 35860 19796 35866 19848
rect 35953 19839 36011 19845
rect 35953 19805 35965 19839
rect 35999 19836 36011 19839
rect 36188 19836 36216 19876
rect 35999 19808 36216 19836
rect 35999 19805 36011 19808
rect 35953 19799 36011 19805
rect 36262 19796 36268 19848
rect 36320 19845 36326 19848
rect 36320 19836 36328 19845
rect 38010 19836 38016 19848
rect 36320 19808 36365 19836
rect 37971 19808 38016 19836
rect 36320 19799 36328 19808
rect 36320 19796 36326 19799
rect 38010 19796 38016 19808
rect 38068 19796 38074 19848
rect 38212 19836 38240 19876
rect 38838 19864 38844 19876
rect 38896 19904 38902 19916
rect 38933 19907 38991 19913
rect 38933 19904 38945 19907
rect 38896 19876 38945 19904
rect 38896 19864 38902 19876
rect 38933 19873 38945 19876
rect 38979 19873 38991 19907
rect 39114 19904 39120 19916
rect 39075 19876 39120 19904
rect 38933 19867 38991 19873
rect 39114 19864 39120 19876
rect 39172 19864 39178 19916
rect 39224 19913 39252 19944
rect 39209 19907 39267 19913
rect 39209 19873 39221 19907
rect 39255 19873 39267 19907
rect 39209 19867 39267 19873
rect 38286 19836 38292 19848
rect 38199 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 39022 19796 39028 19848
rect 39080 19836 39086 19848
rect 39080 19808 39125 19836
rect 39080 19796 39086 19808
rect 34790 19728 34796 19780
rect 34848 19768 34854 19780
rect 36078 19768 36084 19780
rect 34848 19740 36084 19768
rect 34848 19728 34854 19740
rect 36078 19728 36084 19740
rect 36136 19728 36142 19780
rect 36173 19771 36231 19777
rect 36173 19737 36185 19771
rect 36219 19768 36231 19771
rect 37090 19768 37096 19780
rect 36219 19740 37096 19768
rect 36219 19737 36231 19740
rect 36173 19731 36231 19737
rect 37090 19728 37096 19740
rect 37148 19728 37154 19780
rect 38194 19768 38200 19780
rect 38155 19740 38200 19768
rect 38194 19728 38200 19740
rect 38252 19728 38258 19780
rect 36449 19703 36507 19709
rect 36449 19700 36461 19703
rect 34164 19672 36461 19700
rect 36449 19669 36461 19672
rect 36495 19669 36507 19703
rect 36449 19663 36507 19669
rect 39114 19660 39120 19712
rect 39172 19700 39178 19712
rect 48314 19700 48320 19712
rect 39172 19672 48320 19700
rect 39172 19660 39178 19672
rect 48314 19660 48320 19672
rect 48372 19660 48378 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 2041 19499 2099 19505
rect 2041 19465 2053 19499
rect 2087 19496 2099 19499
rect 3789 19499 3847 19505
rect 3789 19496 3801 19499
rect 2087 19468 3801 19496
rect 2087 19465 2099 19468
rect 2041 19459 2099 19465
rect 3789 19465 3801 19468
rect 3835 19465 3847 19499
rect 3789 19459 3847 19465
rect 7193 19499 7251 19505
rect 7193 19465 7205 19499
rect 7239 19496 7251 19499
rect 7239 19468 7696 19496
rect 7239 19465 7251 19468
rect 7193 19459 7251 19465
rect 3697 19431 3755 19437
rect 3697 19397 3709 19431
rect 3743 19428 3755 19431
rect 5166 19428 5172 19440
rect 3743 19400 5172 19428
rect 3743 19397 3755 19400
rect 3697 19391 3755 19397
rect 5166 19388 5172 19400
rect 5224 19388 5230 19440
rect 7668 19437 7696 19468
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7892 19468 8125 19496
rect 7892 19456 7898 19468
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 12805 19499 12863 19505
rect 12805 19465 12817 19499
rect 12851 19465 12863 19499
rect 12805 19459 12863 19465
rect 7653 19431 7711 19437
rect 7653 19397 7665 19431
rect 7699 19397 7711 19431
rect 8202 19428 8208 19440
rect 7653 19391 7711 19397
rect 7852 19400 8208 19428
rect 1394 19320 1400 19372
rect 1452 19360 1458 19372
rect 1581 19363 1639 19369
rect 1581 19360 1593 19363
rect 1452 19332 1593 19360
rect 1452 19320 1458 19332
rect 1581 19329 1593 19332
rect 1627 19329 1639 19363
rect 2222 19360 2228 19372
rect 2183 19332 2228 19360
rect 1581 19323 1639 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 3326 19320 3332 19372
rect 3384 19320 3390 19372
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 6914 19360 6920 19372
rect 6687 19332 6920 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19360 7067 19363
rect 7098 19360 7104 19372
rect 7055 19332 7104 19360
rect 7055 19329 7067 19332
rect 7009 19323 7067 19329
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 7852 19369 7880 19400
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 11790 19428 11796 19440
rect 11532 19400 11796 19428
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8294 19360 8300 19372
rect 7975 19332 8300 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8294 19320 8300 19332
rect 8352 19360 8358 19372
rect 9398 19360 9404 19372
rect 8352 19332 9404 19360
rect 8352 19320 8358 19332
rect 9398 19320 9404 19332
rect 9456 19360 9462 19372
rect 11532 19369 11560 19400
rect 11790 19388 11796 19400
rect 11848 19388 11854 19440
rect 12820 19428 12848 19459
rect 13538 19456 13544 19508
rect 13596 19496 13602 19508
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 13596 19468 15117 19496
rect 13596 19456 13602 19468
rect 15105 19465 15117 19468
rect 15151 19465 15163 19499
rect 15105 19459 15163 19465
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 15930 19496 15936 19508
rect 15436 19468 15936 19496
rect 15436 19456 15442 19468
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 17034 19456 17040 19508
rect 17092 19496 17098 19508
rect 19429 19499 19487 19505
rect 19429 19496 19441 19499
rect 17092 19468 19441 19496
rect 17092 19456 17098 19468
rect 19429 19465 19441 19468
rect 19475 19465 19487 19499
rect 24670 19496 24676 19508
rect 24631 19468 24676 19496
rect 19429 19459 19487 19465
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25038 19496 25044 19508
rect 24999 19468 25044 19496
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 27338 19496 27344 19508
rect 25976 19468 27344 19496
rect 16114 19428 16120 19440
rect 12820 19400 16120 19428
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 17402 19388 17408 19440
rect 17460 19428 17466 19440
rect 20533 19431 20591 19437
rect 20533 19428 20545 19431
rect 17460 19400 20545 19428
rect 17460 19388 17466 19400
rect 20533 19397 20545 19400
rect 20579 19397 20591 19431
rect 25976 19428 26004 19468
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 30561 19499 30619 19505
rect 30561 19465 30573 19499
rect 30607 19496 30619 19499
rect 30742 19496 30748 19508
rect 30607 19468 30748 19496
rect 30607 19465 30619 19468
rect 30561 19459 30619 19465
rect 30742 19456 30748 19468
rect 30800 19456 30806 19508
rect 34054 19496 34060 19508
rect 31036 19468 33548 19496
rect 34015 19468 34060 19496
rect 20533 19391 20591 19397
rect 24872 19400 26004 19428
rect 26053 19431 26111 19437
rect 11517 19363 11575 19369
rect 9456 19332 11468 19360
rect 9456 19320 9462 19332
rect 3344 19233 3372 19320
rect 3878 19292 3884 19304
rect 3839 19264 3884 19292
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 11440 19292 11468 19332
rect 11517 19329 11529 19363
rect 11563 19329 11575 19363
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11517 19323 11575 19329
rect 11624 19332 11713 19360
rect 11624 19292 11652 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 12253 19363 12311 19369
rect 12253 19329 12265 19363
rect 12299 19360 12311 19363
rect 12342 19360 12348 19372
rect 12299 19332 12348 19360
rect 12299 19329 12311 19332
rect 12253 19323 12311 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12952 19332 13277 19360
rect 12952 19320 12958 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13265 19323 13323 19329
rect 11440 19264 11652 19292
rect 3329 19227 3387 19233
rect 3329 19193 3341 19227
rect 3375 19193 3387 19227
rect 8110 19224 8116 19236
rect 3329 19187 3387 19193
rect 7024 19196 8116 19224
rect 7024 19168 7052 19196
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 13280 19224 13308 19323
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13412 19332 13461 19360
rect 13412 19320 13418 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13449 19323 13507 19329
rect 13541 19363 13599 19369
rect 13541 19329 13553 19363
rect 13587 19360 13599 19363
rect 13630 19360 13636 19372
rect 13587 19332 13636 19360
rect 13587 19329 13599 19332
rect 13541 19323 13599 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 15286 19360 15292 19372
rect 15247 19332 15292 19360
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 17126 19360 17132 19372
rect 15519 19332 16436 19360
rect 17087 19332 17132 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 16132 19304 16160 19332
rect 13998 19292 14004 19304
rect 13959 19264 14004 19292
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 13446 19224 13452 19236
rect 13280 19196 13452 19224
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 1397 19159 1455 19165
rect 1397 19125 1409 19159
rect 1443 19156 1455 19159
rect 2682 19156 2688 19168
rect 1443 19128 2688 19156
rect 1443 19125 1455 19128
rect 1397 19119 1455 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 7006 19156 7012 19168
rect 6919 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 7340 19128 7665 19156
rect 7340 19116 7346 19128
rect 7653 19125 7665 19128
rect 7699 19156 7711 19159
rect 8018 19156 8024 19168
rect 7699 19128 8024 19156
rect 7699 19125 7711 19128
rect 7653 19119 7711 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 15396 19156 15424 19255
rect 15580 19224 15608 19255
rect 16114 19252 16120 19304
rect 16172 19252 16178 19304
rect 16408 19292 16436 19332
rect 17126 19320 17132 19332
rect 17184 19320 17190 19372
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18417 19363 18475 19369
rect 18417 19360 18429 19363
rect 18380 19332 18429 19360
rect 18380 19320 18386 19332
rect 18417 19329 18429 19332
rect 18463 19360 18475 19363
rect 19242 19360 19248 19372
rect 18463 19332 19248 19360
rect 18463 19329 18475 19332
rect 18417 19323 18475 19329
rect 19242 19320 19248 19332
rect 19300 19360 19306 19372
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 19300 19332 19809 19360
rect 19300 19320 19306 19332
rect 19797 19329 19809 19332
rect 19843 19360 19855 19363
rect 19843 19332 20668 19360
rect 19843 19329 19855 19332
rect 19797 19323 19855 19329
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 16408 19264 18153 19292
rect 18141 19261 18153 19264
rect 18187 19292 18199 19295
rect 19150 19292 19156 19304
rect 18187 19264 19156 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19518 19252 19524 19304
rect 19576 19292 19582 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19576 19264 19625 19292
rect 19576 19252 19582 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 19702 19252 19708 19304
rect 19760 19292 19766 19304
rect 19760 19264 19805 19292
rect 19760 19252 19766 19264
rect 19886 19252 19892 19304
rect 19944 19292 19950 19304
rect 20640 19292 20668 19332
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 22094 19369 22100 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21692 19332 21833 19360
rect 21692 19320 21698 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22088 19323 22100 19369
rect 22152 19360 22158 19372
rect 24872 19369 24900 19400
rect 26053 19397 26065 19431
rect 26099 19397 26111 19431
rect 26053 19391 26111 19397
rect 24857 19363 24915 19369
rect 22152 19332 22188 19360
rect 22094 19320 22100 19323
rect 22152 19320 22158 19332
rect 24857 19329 24869 19363
rect 24903 19329 24915 19363
rect 25130 19360 25136 19372
rect 25091 19332 25136 19360
rect 24857 19323 24915 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 26068 19334 26096 19391
rect 26234 19388 26240 19440
rect 26292 19437 26298 19440
rect 26292 19431 26311 19437
rect 26299 19397 26311 19431
rect 26292 19391 26311 19397
rect 26973 19431 27031 19437
rect 26973 19397 26985 19431
rect 27019 19397 27031 19431
rect 26973 19391 27031 19397
rect 26292 19388 26298 19391
rect 26988 19360 27016 19391
rect 27154 19388 27160 19440
rect 27212 19437 27218 19440
rect 27212 19431 27231 19437
rect 27219 19397 27231 19431
rect 27212 19391 27231 19397
rect 27212 19388 27218 19391
rect 28718 19388 28724 19440
rect 28776 19428 28782 19440
rect 28776 19400 30420 19428
rect 28776 19388 28782 19400
rect 27982 19360 27988 19372
rect 26068 19306 26188 19334
rect 20898 19292 20904 19304
rect 19944 19264 19989 19292
rect 20640 19264 20904 19292
rect 19944 19252 19950 19264
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 26160 19292 26188 19306
rect 26528 19332 27988 19360
rect 26528 19292 26556 19332
rect 27982 19320 27988 19332
rect 28040 19320 28046 19372
rect 29454 19360 29460 19372
rect 29415 19332 29460 19360
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 29638 19360 29644 19372
rect 29599 19332 29644 19360
rect 29638 19320 29644 19332
rect 29696 19320 29702 19372
rect 30190 19360 30196 19372
rect 30151 19332 30196 19360
rect 30190 19320 30196 19332
rect 30248 19320 30254 19372
rect 30392 19369 30420 19400
rect 30377 19363 30435 19369
rect 30377 19329 30389 19363
rect 30423 19360 30435 19363
rect 30650 19360 30656 19372
rect 30423 19332 30656 19360
rect 30423 19329 30435 19332
rect 30377 19323 30435 19329
rect 30650 19320 30656 19332
rect 30708 19320 30714 19372
rect 26160 19264 26556 19292
rect 28534 19252 28540 19304
rect 28592 19292 28598 19304
rect 30466 19292 30472 19304
rect 28592 19264 30472 19292
rect 28592 19252 28598 19264
rect 30466 19252 30472 19264
rect 30524 19252 30530 19304
rect 30558 19252 30564 19304
rect 30616 19292 30622 19304
rect 31036 19301 31064 19468
rect 31297 19431 31355 19437
rect 31297 19397 31309 19431
rect 31343 19428 31355 19431
rect 31343 19400 32168 19428
rect 31343 19397 31355 19400
rect 31297 19391 31355 19397
rect 31110 19320 31116 19372
rect 31168 19360 31174 19372
rect 31205 19363 31263 19369
rect 31205 19360 31217 19363
rect 31168 19332 31217 19360
rect 31168 19320 31174 19332
rect 31205 19329 31217 19332
rect 31251 19329 31263 19363
rect 31205 19323 31263 19329
rect 31389 19363 31447 19369
rect 31389 19329 31401 19363
rect 31435 19360 31447 19363
rect 32030 19360 32036 19372
rect 31435 19332 32036 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 32030 19320 32036 19332
rect 32088 19320 32094 19372
rect 32140 19369 32168 19400
rect 32125 19363 32183 19369
rect 32125 19329 32137 19363
rect 32171 19360 32183 19363
rect 32582 19360 32588 19372
rect 32171 19332 32588 19360
rect 32171 19329 32183 19332
rect 32125 19323 32183 19329
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 33520 19369 33548 19468
rect 34054 19456 34060 19468
rect 34112 19456 34118 19508
rect 38749 19499 38807 19505
rect 38749 19465 38761 19499
rect 38795 19496 38807 19499
rect 39022 19496 39028 19508
rect 38795 19468 39028 19496
rect 38795 19465 38807 19468
rect 38749 19459 38807 19465
rect 39022 19456 39028 19468
rect 39080 19456 39086 19508
rect 33781 19431 33839 19437
rect 33781 19397 33793 19431
rect 33827 19428 33839 19431
rect 34146 19428 34152 19440
rect 33827 19400 34152 19428
rect 33827 19397 33839 19400
rect 33781 19391 33839 19397
rect 34146 19388 34152 19400
rect 34204 19388 34210 19440
rect 40034 19428 40040 19440
rect 38948 19400 40040 19428
rect 33413 19363 33471 19369
rect 33413 19360 33425 19363
rect 32692 19332 33425 19360
rect 31021 19295 31079 19301
rect 31021 19292 31033 19295
rect 30616 19264 31033 19292
rect 30616 19252 30622 19264
rect 31021 19261 31033 19264
rect 31067 19261 31079 19295
rect 31570 19292 31576 19304
rect 31531 19264 31576 19292
rect 31021 19255 31079 19261
rect 31570 19252 31576 19264
rect 31628 19252 31634 19304
rect 32214 19252 32220 19304
rect 32272 19292 32278 19304
rect 32401 19295 32459 19301
rect 32401 19292 32413 19295
rect 32272 19264 32413 19292
rect 32272 19252 32278 19264
rect 32401 19261 32413 19264
rect 32447 19261 32459 19295
rect 32401 19255 32459 19261
rect 15838 19224 15844 19236
rect 15580 19196 15844 19224
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 20806 19224 20812 19236
rect 16684 19196 20812 19224
rect 16684 19156 16712 19196
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 25498 19184 25504 19236
rect 25556 19224 25562 19236
rect 25777 19227 25835 19233
rect 25777 19224 25789 19227
rect 25556 19196 25789 19224
rect 25556 19184 25562 19196
rect 25777 19193 25789 19196
rect 25823 19224 25835 19227
rect 31938 19224 31944 19236
rect 25823 19196 31944 19224
rect 25823 19193 25835 19196
rect 25777 19187 25835 19193
rect 15396 19128 16712 19156
rect 17221 19159 17279 19165
rect 17221 19125 17233 19159
rect 17267 19156 17279 19159
rect 18046 19156 18052 19168
rect 17267 19128 18052 19156
rect 17267 19125 17279 19128
rect 17221 19119 17279 19125
rect 18046 19116 18052 19128
rect 18104 19156 18110 19168
rect 18414 19156 18420 19168
rect 18104 19128 18420 19156
rect 18104 19116 18110 19128
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 19886 19116 19892 19168
rect 19944 19156 19950 19168
rect 20070 19156 20076 19168
rect 19944 19128 20076 19156
rect 19944 19116 19950 19128
rect 20070 19116 20076 19128
rect 20128 19156 20134 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20128 19128 20637 19156
rect 20128 19116 20134 19128
rect 20625 19125 20637 19128
rect 20671 19156 20683 19159
rect 20990 19156 20996 19168
rect 20671 19128 20996 19156
rect 20671 19125 20683 19128
rect 20625 19119 20683 19125
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 22554 19116 22560 19168
rect 22612 19156 22618 19168
rect 26252 19165 26280 19196
rect 31938 19184 31944 19196
rect 31996 19184 32002 19236
rect 32030 19184 32036 19236
rect 32088 19224 32094 19236
rect 32692 19224 32720 19332
rect 33413 19329 33425 19332
rect 33459 19329 33471 19363
rect 33413 19323 33471 19329
rect 33506 19363 33564 19369
rect 33506 19329 33518 19363
rect 33552 19329 33564 19363
rect 33506 19323 33564 19329
rect 33689 19363 33747 19369
rect 33689 19329 33701 19363
rect 33735 19360 33747 19363
rect 33870 19360 33876 19372
rect 33928 19369 33934 19372
rect 33735 19332 33769 19360
rect 33836 19332 33876 19360
rect 33735 19329 33747 19332
rect 33689 19323 33747 19329
rect 33704 19292 33732 19323
rect 33870 19320 33876 19332
rect 33928 19323 33936 19369
rect 35342 19360 35348 19372
rect 33980 19332 35348 19360
rect 33928 19320 33934 19323
rect 33980 19292 34008 19332
rect 35342 19320 35348 19332
rect 35400 19360 35406 19372
rect 35529 19363 35587 19369
rect 35529 19360 35541 19363
rect 35400 19332 35541 19360
rect 35400 19320 35406 19332
rect 35529 19329 35541 19332
rect 35575 19329 35587 19363
rect 35529 19323 35587 19329
rect 38286 19320 38292 19372
rect 38344 19360 38350 19372
rect 38948 19369 38976 19400
rect 40034 19388 40040 19400
rect 40092 19388 40098 19440
rect 38933 19363 38991 19369
rect 38933 19360 38945 19363
rect 38344 19332 38945 19360
rect 38344 19320 38350 19332
rect 38933 19329 38945 19332
rect 38979 19329 38991 19363
rect 38933 19323 38991 19329
rect 39117 19363 39175 19369
rect 39117 19329 39129 19363
rect 39163 19329 39175 19363
rect 39117 19323 39175 19329
rect 39209 19363 39267 19369
rect 39209 19329 39221 19363
rect 39255 19329 39267 19363
rect 39209 19323 39267 19329
rect 33704 19264 34008 19292
rect 34790 19252 34796 19304
rect 34848 19292 34854 19304
rect 35253 19295 35311 19301
rect 35253 19292 35265 19295
rect 34848 19264 35265 19292
rect 34848 19252 34854 19264
rect 35253 19261 35265 19264
rect 35299 19261 35311 19295
rect 35253 19255 35311 19261
rect 38194 19252 38200 19304
rect 38252 19292 38258 19304
rect 39132 19292 39160 19323
rect 38252 19264 39160 19292
rect 38252 19252 38258 19264
rect 32088 19196 32720 19224
rect 32088 19184 32094 19196
rect 38010 19184 38016 19236
rect 38068 19224 38074 19236
rect 39224 19224 39252 19323
rect 38068 19196 39252 19224
rect 38068 19184 38074 19196
rect 23201 19159 23259 19165
rect 23201 19156 23213 19159
rect 22612 19128 23213 19156
rect 22612 19116 22618 19128
rect 23201 19125 23213 19128
rect 23247 19125 23259 19159
rect 23201 19119 23259 19125
rect 26237 19159 26295 19165
rect 26237 19125 26249 19159
rect 26283 19125 26295 19159
rect 26418 19156 26424 19168
rect 26379 19128 26424 19156
rect 26237 19119 26295 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 27062 19116 27068 19168
rect 27120 19156 27126 19168
rect 27157 19159 27215 19165
rect 27157 19156 27169 19159
rect 27120 19128 27169 19156
rect 27120 19116 27126 19128
rect 27157 19125 27169 19128
rect 27203 19156 27215 19159
rect 27709 19159 27767 19165
rect 27709 19156 27721 19159
rect 27203 19128 27721 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 27709 19125 27721 19128
rect 27755 19156 27767 19159
rect 29362 19156 29368 19168
rect 27755 19128 29368 19156
rect 27755 19125 27767 19128
rect 27709 19119 27767 19125
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 29549 19159 29607 19165
rect 29549 19125 29561 19159
rect 29595 19156 29607 19159
rect 30006 19156 30012 19168
rect 29595 19128 30012 19156
rect 29595 19125 29607 19128
rect 29549 19119 29607 19125
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 36078 19116 36084 19168
rect 36136 19156 36142 19168
rect 36998 19156 37004 19168
rect 36136 19128 37004 19156
rect 36136 19116 36142 19128
rect 36998 19116 37004 19128
rect 37056 19116 37062 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 3142 18952 3148 18964
rect 3055 18924 3148 18952
rect 3142 18912 3148 18924
rect 3200 18952 3206 18964
rect 7006 18952 7012 18964
rect 3200 18924 7012 18952
rect 3200 18912 3206 18924
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 7374 18952 7380 18964
rect 7239 18924 7380 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 10413 18955 10471 18961
rect 10413 18921 10425 18955
rect 10459 18952 10471 18955
rect 17126 18952 17132 18964
rect 10459 18924 17132 18952
rect 10459 18921 10471 18924
rect 10413 18915 10471 18921
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 19518 18952 19524 18964
rect 19479 18924 19524 18952
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 19886 18952 19892 18964
rect 19628 18924 19892 18952
rect 7742 18884 7748 18896
rect 6840 18856 7748 18884
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 6840 18757 6868 18856
rect 7742 18844 7748 18856
rect 7800 18884 7806 18896
rect 11977 18887 12035 18893
rect 7800 18856 10548 18884
rect 7800 18844 7806 18856
rect 6914 18776 6920 18828
rect 6972 18816 6978 18828
rect 7101 18819 7159 18825
rect 7101 18816 7113 18819
rect 6972 18788 7113 18816
rect 6972 18776 6978 18788
rect 7101 18785 7113 18788
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 8904 18788 9168 18816
rect 8904 18776 8910 18788
rect 1765 18751 1823 18757
rect 1765 18748 1777 18751
rect 1544 18720 1777 18748
rect 1544 18708 1550 18720
rect 1765 18717 1777 18720
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 7837 18751 7895 18757
rect 7837 18748 7849 18751
rect 7432 18720 7849 18748
rect 7432 18708 7438 18720
rect 7837 18717 7849 18720
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7984 18720 8033 18748
rect 7984 18708 7990 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9140 18757 9168 18788
rect 10520 18757 10548 18856
rect 11977 18853 11989 18887
rect 12023 18884 12035 18887
rect 12526 18884 12532 18896
rect 12023 18856 12532 18884
rect 12023 18853 12035 18856
rect 11977 18847 12035 18853
rect 12526 18844 12532 18856
rect 12584 18884 12590 18896
rect 15838 18884 15844 18896
rect 12584 18856 15844 18884
rect 12584 18844 12590 18856
rect 15838 18844 15844 18856
rect 15896 18884 15902 18896
rect 17034 18884 17040 18896
rect 15896 18856 17040 18884
rect 15896 18844 15902 18856
rect 17034 18844 17040 18856
rect 17092 18844 17098 18896
rect 17144 18816 17172 18912
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 19628 18884 19656 18924
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 20530 18952 20536 18964
rect 20491 18924 20536 18952
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22189 18955 22247 18961
rect 22189 18952 22201 18955
rect 22152 18924 22201 18952
rect 22152 18912 22158 18924
rect 22189 18921 22201 18924
rect 22235 18921 22247 18955
rect 22189 18915 22247 18921
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 28718 18952 28724 18964
rect 22428 18924 28724 18952
rect 22428 18912 22434 18924
rect 28718 18912 28724 18924
rect 28776 18912 28782 18964
rect 28810 18912 28816 18964
rect 28868 18952 28874 18964
rect 28994 18952 29000 18964
rect 28868 18924 28913 18952
rect 28955 18924 29000 18952
rect 28868 18912 28874 18924
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 29549 18955 29607 18961
rect 29549 18921 29561 18955
rect 29595 18952 29607 18955
rect 30190 18952 30196 18964
rect 29595 18924 30196 18952
rect 29595 18921 29607 18924
rect 29549 18915 29607 18921
rect 30190 18912 30196 18924
rect 30248 18912 30254 18964
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 36630 18952 36636 18964
rect 30524 18924 36636 18952
rect 30524 18912 30530 18924
rect 36630 18912 36636 18924
rect 36688 18912 36694 18964
rect 18012 18856 19656 18884
rect 18012 18844 18018 18856
rect 25130 18844 25136 18896
rect 25188 18884 25194 18896
rect 25406 18884 25412 18896
rect 25188 18856 25412 18884
rect 25188 18844 25194 18856
rect 25406 18844 25412 18856
rect 25464 18844 25470 18896
rect 28902 18844 28908 18896
rect 28960 18884 28966 18896
rect 32677 18887 32735 18893
rect 32677 18884 32689 18887
rect 28960 18856 32689 18884
rect 28960 18844 28966 18856
rect 32677 18853 32689 18856
rect 32723 18853 32735 18887
rect 36170 18884 36176 18896
rect 32677 18847 32735 18853
rect 34992 18856 36176 18884
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 11808 18788 14136 18816
rect 17144 18788 17417 18816
rect 11808 18757 11836 18788
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8720 18720 8953 18748
rect 8720 18708 8726 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 11793 18711 11851 18717
rect 2032 18683 2090 18689
rect 2032 18649 2044 18683
rect 2078 18680 2090 18683
rect 3786 18680 3792 18692
rect 2078 18652 3792 18680
rect 2078 18649 2090 18652
rect 2032 18643 2090 18649
rect 3786 18640 3792 18652
rect 3844 18640 3850 18692
rect 8202 18680 8208 18692
rect 8163 18652 8208 18680
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 9033 18683 9091 18689
rect 9033 18649 9045 18683
rect 9079 18680 9091 18683
rect 10336 18680 10364 18711
rect 10686 18680 10692 18692
rect 9079 18652 10692 18680
rect 9079 18649 9091 18652
rect 9033 18643 9091 18649
rect 10686 18640 10692 18652
rect 10744 18640 10750 18692
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 6822 18612 6828 18624
rect 1820 18584 6828 18612
rect 1820 18572 1826 18584
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 7377 18615 7435 18621
rect 7377 18612 7389 18615
rect 6972 18584 7389 18612
rect 6972 18572 6978 18584
rect 7377 18581 7389 18584
rect 7423 18581 7435 18615
rect 7377 18575 7435 18581
rect 10226 18572 10232 18624
rect 10284 18612 10290 18624
rect 11808 18612 11836 18711
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 14108 18757 14136 18788
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 18598 18816 18604 18828
rect 17727 18788 18604 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 18598 18776 18604 18788
rect 18656 18816 18662 18828
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 18656 18788 19993 18816
rect 18656 18776 18662 18788
rect 19981 18785 19993 18788
rect 20027 18816 20039 18819
rect 20254 18816 20260 18828
rect 20027 18788 20260 18816
rect 20027 18785 20039 18788
rect 19981 18779 20039 18785
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 20809 18819 20867 18825
rect 20809 18785 20821 18819
rect 20855 18816 20867 18819
rect 22186 18816 22192 18828
rect 20855 18788 22192 18816
rect 20855 18785 20867 18788
rect 20809 18779 20867 18785
rect 22186 18776 22192 18788
rect 22244 18776 22250 18828
rect 22554 18816 22560 18828
rect 22296 18788 22560 18816
rect 14093 18751 14151 18757
rect 14093 18717 14105 18751
rect 14139 18748 14151 18751
rect 17310 18748 17316 18760
rect 14139 18720 17316 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 19702 18748 19708 18760
rect 19663 18720 19708 18748
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 19797 18751 19855 18757
rect 19797 18717 19809 18751
rect 19843 18717 19855 18751
rect 19797 18711 19855 18717
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 20714 18748 20720 18760
rect 20675 18720 20720 18748
rect 19889 18711 19947 18717
rect 15562 18680 15568 18692
rect 15475 18652 15568 18680
rect 15562 18640 15568 18652
rect 15620 18680 15626 18692
rect 15620 18652 16712 18680
rect 15620 18640 15626 18652
rect 12710 18612 12716 18624
rect 10284 18584 11836 18612
rect 12623 18584 12716 18612
rect 10284 18572 10290 18584
rect 12710 18572 12716 18584
rect 12768 18612 12774 18624
rect 12894 18612 12900 18624
rect 12768 18584 12900 18612
rect 12768 18572 12774 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14277 18615 14335 18621
rect 14277 18581 14289 18615
rect 14323 18612 14335 18615
rect 15746 18612 15752 18624
rect 14323 18584 15752 18612
rect 14323 18581 14335 18584
rect 14277 18575 14335 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 15841 18615 15899 18621
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 15930 18612 15936 18624
rect 15887 18584 15936 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 16684 18612 16712 18652
rect 19242 18640 19248 18692
rect 19300 18680 19306 18692
rect 19812 18680 19840 18711
rect 19300 18652 19840 18680
rect 19904 18680 19932 18711
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 20898 18748 20904 18760
rect 20859 18720 20904 18748
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21048 18720 21093 18748
rect 21048 18708 21054 18720
rect 22296 18680 22324 18788
rect 22554 18776 22560 18788
rect 22612 18776 22618 18828
rect 25148 18816 25176 18844
rect 22664 18788 25176 18816
rect 22664 18760 22692 18788
rect 30098 18776 30104 18828
rect 30156 18816 30162 18828
rect 30156 18788 30236 18816
rect 30156 18776 30162 18788
rect 22370 18708 22376 18760
rect 22428 18748 22434 18760
rect 22646 18748 22652 18760
rect 22428 18720 22473 18748
rect 22559 18720 22652 18748
rect 22428 18708 22434 18720
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 22756 18720 28764 18748
rect 22756 18680 22784 18720
rect 19904 18652 22324 18680
rect 22480 18652 22784 18680
rect 19300 18640 19306 18652
rect 22480 18612 22508 18652
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25225 18683 25283 18689
rect 25225 18680 25237 18683
rect 25188 18652 25237 18680
rect 25188 18640 25194 18652
rect 25225 18649 25237 18652
rect 25271 18680 25283 18683
rect 26142 18680 26148 18692
rect 25271 18652 26148 18680
rect 25271 18649 25283 18652
rect 25225 18643 25283 18649
rect 26142 18640 26148 18652
rect 26200 18640 26206 18692
rect 28626 18680 28632 18692
rect 28587 18652 28632 18680
rect 28626 18640 28632 18652
rect 28684 18640 28690 18692
rect 28736 18680 28764 18720
rect 29178 18708 29184 18760
rect 29236 18748 29242 18760
rect 29805 18751 29863 18757
rect 29805 18748 29817 18751
rect 29236 18720 29817 18748
rect 29236 18708 29242 18720
rect 29805 18717 29817 18720
rect 29851 18717 29863 18751
rect 29805 18711 29863 18717
rect 29914 18748 29972 18754
rect 29914 18714 29926 18748
rect 29960 18714 29972 18748
rect 29914 18708 29972 18714
rect 30006 18708 30012 18760
rect 30064 18757 30070 18760
rect 30208 18757 30236 18788
rect 31846 18776 31852 18828
rect 31904 18816 31910 18828
rect 31904 18788 32352 18816
rect 31904 18776 31910 18788
rect 30064 18748 30072 18757
rect 30193 18751 30251 18757
rect 30064 18720 30109 18748
rect 30064 18711 30072 18720
rect 30193 18717 30205 18751
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 30064 18708 30070 18711
rect 30926 18708 30932 18760
rect 30984 18748 30990 18760
rect 32030 18748 32036 18760
rect 30984 18720 32036 18748
rect 30984 18708 30990 18720
rect 32030 18708 32036 18720
rect 32088 18708 32094 18760
rect 32214 18757 32220 18760
rect 32181 18751 32220 18757
rect 32181 18717 32193 18751
rect 32181 18711 32220 18717
rect 32214 18708 32220 18711
rect 32272 18708 32278 18760
rect 32324 18757 32352 18788
rect 33502 18776 33508 18828
rect 33560 18816 33566 18828
rect 34992 18825 35020 18856
rect 36170 18844 36176 18856
rect 36228 18844 36234 18896
rect 38654 18884 38660 18896
rect 36372 18856 38660 18884
rect 34701 18819 34759 18825
rect 34701 18816 34713 18819
rect 33560 18788 34713 18816
rect 33560 18776 33566 18788
rect 34701 18785 34713 18788
rect 34747 18785 34759 18819
rect 34701 18779 34759 18785
rect 34977 18819 35035 18825
rect 34977 18785 34989 18819
rect 35023 18785 35035 18819
rect 36372 18816 36400 18856
rect 38654 18844 38660 18856
rect 38712 18884 38718 18896
rect 39853 18887 39911 18893
rect 39853 18884 39865 18887
rect 38712 18856 39865 18884
rect 38712 18844 38718 18856
rect 39853 18853 39865 18856
rect 39899 18853 39911 18887
rect 39853 18847 39911 18853
rect 34977 18779 35035 18785
rect 36152 18788 36400 18816
rect 36648 18788 37693 18816
rect 32309 18751 32367 18757
rect 32309 18717 32321 18751
rect 32355 18717 32367 18751
rect 32309 18711 32367 18717
rect 32539 18751 32597 18757
rect 32539 18717 32551 18751
rect 32585 18748 32597 18751
rect 32766 18748 32772 18760
rect 32585 18720 32772 18748
rect 32585 18717 32597 18720
rect 32539 18711 32597 18717
rect 32766 18708 32772 18720
rect 32824 18748 32830 18760
rect 33870 18748 33876 18760
rect 32824 18720 33876 18748
rect 32824 18708 32830 18720
rect 33870 18708 33876 18720
rect 33928 18708 33934 18760
rect 35986 18748 35992 18760
rect 35947 18720 35992 18748
rect 35986 18708 35992 18720
rect 36044 18708 36050 18760
rect 36152 18757 36180 18788
rect 36648 18760 36676 18788
rect 36137 18751 36195 18757
rect 36137 18717 36149 18751
rect 36183 18717 36195 18751
rect 36137 18711 36195 18717
rect 36495 18751 36553 18757
rect 36495 18717 36507 18751
rect 36541 18748 36553 18751
rect 36630 18748 36636 18760
rect 36541 18720 36636 18748
rect 36541 18717 36553 18720
rect 36495 18711 36553 18717
rect 36630 18708 36636 18720
rect 36688 18708 36694 18760
rect 37182 18748 37188 18760
rect 37143 18720 37188 18748
rect 37182 18708 37188 18720
rect 37240 18708 37246 18760
rect 37366 18757 37372 18760
rect 37333 18751 37372 18757
rect 37333 18717 37345 18751
rect 37333 18711 37372 18717
rect 37366 18708 37372 18711
rect 37424 18708 37430 18760
rect 37665 18757 37693 18788
rect 37650 18751 37708 18757
rect 37650 18717 37662 18751
rect 37696 18717 37708 18751
rect 40034 18748 40040 18760
rect 39995 18720 40040 18748
rect 37650 18711 37708 18717
rect 40034 18708 40040 18720
rect 40092 18708 40098 18760
rect 29546 18680 29552 18692
rect 28736 18652 29552 18680
rect 29546 18640 29552 18652
rect 29604 18640 29610 18692
rect 16684 18584 22508 18612
rect 22554 18572 22560 18624
rect 22612 18612 22618 18624
rect 22612 18584 22657 18612
rect 22612 18572 22618 18584
rect 24394 18572 24400 18624
rect 24452 18612 24458 18624
rect 27062 18612 27068 18624
rect 24452 18584 27068 18612
rect 24452 18572 24458 18584
rect 27062 18572 27068 18584
rect 27120 18612 27126 18624
rect 27890 18612 27896 18624
rect 27120 18584 27896 18612
rect 27120 18572 27126 18584
rect 27890 18572 27896 18584
rect 27948 18572 27954 18624
rect 28839 18615 28897 18621
rect 28839 18581 28851 18615
rect 28885 18612 28897 18615
rect 29454 18612 29460 18624
rect 28885 18584 29460 18612
rect 28885 18581 28897 18584
rect 28839 18575 28897 18581
rect 29454 18572 29460 18584
rect 29512 18612 29518 18624
rect 29929 18612 29957 18708
rect 32401 18683 32459 18689
rect 32401 18649 32413 18683
rect 32447 18680 32459 18683
rect 36265 18683 36323 18689
rect 36265 18680 36277 18683
rect 32447 18652 32628 18680
rect 32447 18649 32459 18652
rect 32401 18643 32459 18649
rect 32600 18624 32628 18652
rect 36096 18652 36277 18680
rect 36096 18624 36124 18652
rect 36265 18649 36277 18652
rect 36311 18649 36323 18683
rect 36265 18643 36323 18649
rect 36357 18683 36415 18689
rect 36357 18649 36369 18683
rect 36403 18680 36415 18683
rect 36906 18680 36912 18692
rect 36403 18652 36912 18680
rect 36403 18649 36415 18652
rect 36357 18643 36415 18649
rect 36906 18640 36912 18652
rect 36964 18640 36970 18692
rect 36998 18640 37004 18692
rect 37056 18680 37062 18692
rect 37461 18683 37519 18689
rect 37461 18680 37473 18683
rect 37056 18652 37473 18680
rect 37056 18640 37062 18652
rect 37461 18649 37473 18652
rect 37507 18649 37519 18683
rect 37461 18643 37519 18649
rect 37550 18640 37556 18692
rect 37608 18680 37614 18692
rect 37608 18652 37653 18680
rect 37608 18640 37614 18652
rect 39942 18640 39948 18692
rect 40000 18680 40006 18692
rect 40129 18683 40187 18689
rect 40129 18680 40141 18683
rect 40000 18652 40141 18680
rect 40000 18640 40006 18652
rect 40129 18649 40141 18652
rect 40175 18649 40187 18683
rect 40129 18643 40187 18649
rect 29512 18584 29957 18612
rect 29512 18572 29518 18584
rect 32582 18572 32588 18624
rect 32640 18572 32646 18624
rect 36078 18572 36084 18624
rect 36136 18572 36142 18624
rect 36630 18612 36636 18624
rect 36591 18584 36636 18612
rect 36630 18572 36636 18584
rect 36688 18572 36694 18624
rect 37826 18612 37832 18624
rect 37787 18584 37832 18612
rect 37826 18572 37832 18584
rect 37884 18572 37890 18624
rect 38010 18572 38016 18624
rect 38068 18612 38074 18624
rect 40221 18615 40279 18621
rect 40221 18612 40233 18615
rect 38068 18584 40233 18612
rect 38068 18572 38074 18584
rect 40221 18581 40233 18584
rect 40267 18581 40279 18615
rect 40402 18612 40408 18624
rect 40363 18584 40408 18612
rect 40221 18575 40279 18581
rect 40402 18572 40408 18584
rect 40460 18572 40466 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 2593 18411 2651 18417
rect 2593 18377 2605 18411
rect 2639 18408 2651 18411
rect 3142 18408 3148 18420
rect 2639 18380 3148 18408
rect 2639 18377 2651 18380
rect 2593 18371 2651 18377
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 3878 18408 3884 18420
rect 3839 18380 3884 18408
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 9674 18408 9680 18420
rect 9635 18380 9680 18408
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 15562 18408 15568 18420
rect 11931 18380 15568 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 18322 18408 18328 18420
rect 17276 18380 18328 18408
rect 17276 18368 17282 18380
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20714 18408 20720 18420
rect 20027 18380 20720 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 37826 18408 37832 18420
rect 20864 18380 37832 18408
rect 20864 18368 20870 18380
rect 37826 18368 37832 18380
rect 37884 18368 37890 18420
rect 2682 18340 2688 18352
rect 2643 18312 2688 18340
rect 2682 18300 2688 18312
rect 2740 18300 2746 18352
rect 10134 18340 10140 18352
rect 8312 18312 10140 18340
rect 1397 18275 1455 18281
rect 1397 18241 1409 18275
rect 1443 18241 1455 18275
rect 1397 18235 1455 18241
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 4614 18272 4620 18284
rect 3835 18244 4620 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 1412 18136 1440 18235
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 6914 18272 6920 18284
rect 6875 18244 6920 18272
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7834 18232 7840 18284
rect 7892 18272 7898 18284
rect 8312 18281 8340 18312
rect 10134 18300 10140 18312
rect 10192 18300 10198 18352
rect 15746 18300 15752 18352
rect 15804 18340 15810 18352
rect 22370 18340 22376 18352
rect 15804 18312 17356 18340
rect 15804 18300 15810 18312
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 7892 18244 8309 18272
rect 7892 18232 7898 18244
rect 8297 18241 8309 18244
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 8564 18275 8622 18281
rect 8564 18241 8576 18275
rect 8610 18272 8622 18275
rect 8938 18272 8944 18284
rect 8610 18244 8944 18272
rect 8610 18241 8622 18244
rect 8564 18235 8622 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18272 11759 18275
rect 12342 18272 12348 18284
rect 11747 18244 12348 18272
rect 11747 18241 11759 18244
rect 11701 18235 11759 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 15470 18272 15476 18284
rect 15431 18244 15476 18272
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16114 18272 16120 18284
rect 15703 18244 16120 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16114 18232 16120 18244
rect 16172 18272 16178 18284
rect 16666 18272 16672 18284
rect 16172 18244 16672 18272
rect 16172 18232 16178 18244
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 17218 18272 17224 18284
rect 17179 18244 17224 18272
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17328 18272 17356 18312
rect 18616 18312 19472 18340
rect 18616 18284 18644 18312
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 17328 18244 18245 18272
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 18598 18272 18604 18284
rect 18371 18244 18604 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19444 18281 19472 18312
rect 19904 18312 22376 18340
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19116 18244 19165 18272
rect 19116 18232 19122 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19430 18275 19488 18281
rect 19430 18241 19442 18275
rect 19476 18241 19488 18275
rect 19430 18235 19488 18241
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3050 18204 3056 18216
rect 2915 18176 3056 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3050 18164 3056 18176
rect 3108 18204 3114 18216
rect 3878 18204 3884 18216
rect 3108 18176 3884 18204
rect 3108 18164 3114 18176
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 11422 18164 11428 18216
rect 11480 18204 11486 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 11480 18176 11529 18204
rect 11480 18164 11486 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 15194 18164 15200 18216
rect 15252 18204 15258 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 15252 18176 16865 18204
rect 15252 18164 15258 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 6178 18136 6184 18148
rect 1412 18108 6184 18136
rect 6178 18096 6184 18108
rect 6236 18096 6242 18148
rect 14458 18096 14464 18148
rect 14516 18136 14522 18148
rect 17052 18136 17080 18167
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17313 18207 17371 18213
rect 17184 18176 17229 18204
rect 17184 18164 17190 18176
rect 17313 18173 17325 18207
rect 17359 18204 17371 18207
rect 17954 18204 17960 18216
rect 17359 18176 17960 18204
rect 17359 18173 17371 18176
rect 17313 18167 17371 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 17865 18139 17923 18145
rect 17865 18136 17877 18139
rect 14516 18108 16988 18136
rect 17052 18108 17877 18136
rect 14516 18096 14522 18108
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 3326 18068 3332 18080
rect 2271 18040 3332 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 7101 18071 7159 18077
rect 7101 18037 7113 18071
rect 7147 18068 7159 18071
rect 8018 18068 8024 18080
rect 7147 18040 8024 18068
rect 7147 18037 7159 18040
rect 7101 18031 7159 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 16960 18068 16988 18108
rect 17865 18105 17877 18108
rect 17911 18105 17923 18139
rect 18064 18136 18092 18167
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 19242 18204 19248 18216
rect 18196 18176 19248 18204
rect 18196 18164 18202 18176
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19904 18204 19932 18312
rect 22370 18300 22376 18312
rect 22428 18300 22434 18352
rect 30834 18340 30840 18352
rect 26896 18312 30840 18340
rect 19978 18232 19984 18284
rect 20036 18272 20042 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20036 18244 20177 18272
rect 20036 18232 20042 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18272 20407 18275
rect 22002 18272 22008 18284
rect 20395 18244 22008 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 19383 18176 19932 18204
rect 20257 18207 20315 18213
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 20438 18204 20444 18216
rect 20399 18176 20444 18204
rect 20257 18167 20315 18173
rect 19058 18136 19064 18148
rect 18064 18108 19064 18136
rect 17865 18099 17923 18105
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19260 18136 19288 18164
rect 20272 18136 20300 18167
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 20622 18164 20628 18216
rect 20680 18204 20686 18216
rect 26896 18204 26924 18312
rect 30834 18300 30840 18312
rect 30892 18300 30898 18352
rect 31202 18340 31208 18352
rect 31163 18312 31208 18340
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 31297 18343 31355 18349
rect 31297 18309 31309 18343
rect 31343 18340 31355 18343
rect 31570 18340 31576 18352
rect 31343 18312 31576 18340
rect 31343 18309 31355 18312
rect 31297 18303 31355 18309
rect 31570 18300 31576 18312
rect 31628 18300 31634 18352
rect 37366 18300 37372 18352
rect 37424 18340 37430 18352
rect 38841 18343 38899 18349
rect 37424 18312 38792 18340
rect 37424 18300 37430 18312
rect 27062 18272 27068 18284
rect 27023 18244 27068 18272
rect 27062 18232 27068 18244
rect 27120 18232 27126 18284
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27321 18275 27379 18281
rect 27321 18272 27333 18275
rect 27212 18244 27333 18272
rect 27212 18232 27218 18244
rect 27321 18241 27333 18244
rect 27367 18241 27379 18275
rect 27321 18235 27379 18241
rect 28997 18275 29055 18281
rect 28997 18241 29009 18275
rect 29043 18272 29055 18275
rect 29178 18272 29184 18284
rect 29043 18244 29077 18272
rect 29139 18244 29184 18272
rect 29043 18241 29055 18244
rect 28997 18235 29055 18241
rect 28626 18204 28632 18216
rect 20680 18176 26924 18204
rect 28460 18176 28632 18204
rect 20680 18164 20686 18176
rect 22278 18136 22284 18148
rect 19260 18108 20300 18136
rect 22066 18108 22284 18136
rect 18138 18068 18144 18080
rect 16960 18040 18144 18068
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18969 18071 19027 18077
rect 18969 18068 18981 18071
rect 18380 18040 18981 18068
rect 18380 18028 18386 18040
rect 18969 18037 18981 18040
rect 19015 18037 19027 18071
rect 18969 18031 19027 18037
rect 21542 18028 21548 18080
rect 21600 18068 21606 18080
rect 22066 18068 22094 18108
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 28460 18145 28488 18176
rect 28626 18164 28632 18176
rect 28684 18204 28690 18216
rect 29012 18204 29040 18235
rect 29178 18232 29184 18244
rect 29236 18232 29242 18284
rect 29273 18275 29331 18281
rect 29273 18241 29285 18275
rect 29319 18272 29331 18275
rect 29454 18272 29460 18284
rect 29319 18244 29460 18272
rect 29319 18241 29331 18244
rect 29273 18235 29331 18241
rect 29454 18232 29460 18244
rect 29512 18272 29518 18284
rect 30374 18272 30380 18284
rect 29512 18244 30380 18272
rect 29512 18232 29518 18244
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 30926 18272 30932 18284
rect 30887 18244 30932 18272
rect 30926 18232 30932 18244
rect 30984 18232 30990 18284
rect 31110 18281 31116 18284
rect 31077 18275 31116 18281
rect 31077 18241 31089 18275
rect 31077 18235 31116 18241
rect 31092 18232 31116 18235
rect 31168 18232 31174 18284
rect 31435 18275 31493 18281
rect 31435 18241 31447 18275
rect 31481 18272 31493 18275
rect 31662 18272 31668 18284
rect 31481 18244 31668 18272
rect 31481 18241 31493 18244
rect 31435 18235 31493 18241
rect 31662 18232 31668 18244
rect 31720 18232 31726 18284
rect 33502 18232 33508 18284
rect 33560 18272 33566 18284
rect 33597 18275 33655 18281
rect 33597 18272 33609 18275
rect 33560 18244 33609 18272
rect 33560 18232 33566 18244
rect 33597 18241 33609 18244
rect 33643 18241 33655 18275
rect 33597 18235 33655 18241
rect 35161 18275 35219 18281
rect 35161 18241 35173 18275
rect 35207 18272 35219 18275
rect 35802 18272 35808 18284
rect 35207 18244 35808 18272
rect 35207 18241 35219 18244
rect 35161 18235 35219 18241
rect 35802 18232 35808 18244
rect 35860 18232 35866 18284
rect 35986 18232 35992 18284
rect 36044 18272 36050 18284
rect 37182 18272 37188 18284
rect 36044 18244 37188 18272
rect 36044 18232 36050 18244
rect 37182 18232 37188 18244
rect 37240 18232 37246 18284
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18272 37335 18275
rect 37323 18244 37412 18272
rect 37323 18241 37335 18244
rect 37277 18235 37335 18241
rect 31092 18204 31120 18232
rect 28684 18176 31120 18204
rect 28684 18164 28690 18176
rect 32122 18164 32128 18216
rect 32180 18204 32186 18216
rect 32309 18207 32367 18213
rect 32309 18204 32321 18207
rect 32180 18176 32321 18204
rect 32180 18164 32186 18176
rect 32309 18173 32321 18176
rect 32355 18173 32367 18207
rect 32309 18167 32367 18173
rect 32585 18207 32643 18213
rect 32585 18173 32597 18207
rect 32631 18173 32643 18207
rect 33870 18204 33876 18216
rect 33831 18176 33876 18204
rect 32585 18167 32643 18173
rect 28445 18139 28503 18145
rect 28445 18105 28457 18139
rect 28491 18105 28503 18139
rect 30282 18136 30288 18148
rect 28445 18099 28503 18105
rect 28552 18108 30288 18136
rect 21600 18040 22094 18068
rect 21600 18028 21606 18040
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 28552 18068 28580 18108
rect 30282 18096 30288 18108
rect 30340 18096 30346 18148
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 32600 18136 32628 18167
rect 33870 18164 33876 18176
rect 33928 18164 33934 18216
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 34885 18207 34943 18213
rect 34885 18204 34897 18207
rect 34848 18176 34897 18204
rect 34848 18164 34854 18176
rect 34885 18173 34897 18176
rect 34931 18173 34943 18207
rect 37384 18204 37412 18244
rect 37458 18232 37464 18284
rect 37516 18272 37522 18284
rect 38764 18272 38792 18312
rect 38841 18309 38853 18343
rect 38887 18340 38899 18343
rect 38930 18340 38936 18352
rect 38887 18312 38936 18340
rect 38887 18309 38899 18312
rect 38841 18303 38899 18309
rect 38930 18300 38936 18312
rect 38988 18340 38994 18352
rect 39942 18340 39948 18352
rect 38988 18312 39948 18340
rect 38988 18300 38994 18312
rect 39942 18300 39948 18312
rect 40000 18300 40006 18352
rect 39669 18275 39727 18281
rect 39669 18272 39681 18275
rect 37516 18244 38240 18272
rect 38764 18244 39681 18272
rect 37516 18232 37522 18244
rect 38212 18216 38240 18244
rect 39669 18241 39681 18244
rect 39715 18241 39727 18275
rect 39669 18235 39727 18241
rect 38010 18204 38016 18216
rect 37384 18176 38016 18204
rect 34885 18167 34943 18173
rect 38010 18164 38016 18176
rect 38068 18164 38074 18216
rect 38194 18164 38200 18216
rect 38252 18204 38258 18216
rect 39025 18207 39083 18213
rect 39025 18204 39037 18207
rect 38252 18176 39037 18204
rect 38252 18164 38258 18176
rect 39025 18173 39037 18176
rect 39071 18173 39083 18207
rect 39025 18167 39083 18173
rect 33962 18136 33968 18148
rect 30432 18108 33968 18136
rect 30432 18096 30438 18108
rect 33962 18096 33968 18108
rect 34020 18096 34026 18148
rect 39684 18136 39712 18235
rect 40034 18232 40040 18284
rect 40092 18272 40098 18284
rect 40753 18275 40811 18281
rect 40753 18272 40765 18275
rect 40092 18244 40765 18272
rect 40092 18232 40098 18244
rect 40753 18241 40765 18244
rect 40799 18241 40811 18275
rect 40753 18235 40811 18241
rect 39761 18207 39819 18213
rect 39761 18173 39773 18207
rect 39807 18204 39819 18207
rect 40402 18204 40408 18216
rect 39807 18176 40408 18204
rect 39807 18173 39819 18176
rect 39761 18167 39819 18173
rect 40402 18164 40408 18176
rect 40460 18164 40466 18216
rect 40494 18164 40500 18216
rect 40552 18204 40558 18216
rect 40552 18176 40597 18204
rect 40552 18164 40558 18176
rect 39684 18108 40448 18136
rect 22244 18040 28580 18068
rect 28997 18071 29055 18077
rect 22244 18028 22250 18040
rect 28997 18037 29009 18071
rect 29043 18068 29055 18071
rect 29546 18068 29552 18080
rect 29043 18040 29552 18068
rect 29043 18037 29055 18040
rect 28997 18031 29055 18037
rect 29546 18028 29552 18040
rect 29604 18028 29610 18080
rect 31478 18028 31484 18080
rect 31536 18068 31542 18080
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 31536 18040 31585 18068
rect 31536 18028 31542 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 37366 18068 37372 18080
rect 37327 18040 37372 18068
rect 31573 18031 31631 18037
rect 37366 18028 37372 18040
rect 37424 18028 37430 18080
rect 40037 18071 40095 18077
rect 40037 18037 40049 18071
rect 40083 18068 40095 18071
rect 40310 18068 40316 18080
rect 40083 18040 40316 18068
rect 40083 18037 40095 18040
rect 40037 18031 40095 18037
rect 40310 18028 40316 18040
rect 40368 18028 40374 18080
rect 40420 18068 40448 18108
rect 41877 18071 41935 18077
rect 41877 18068 41889 18071
rect 40420 18040 41889 18068
rect 41877 18037 41889 18040
rect 41923 18037 41935 18071
rect 41877 18031 41935 18037
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 6178 17864 6184 17876
rect 2746 17836 5764 17864
rect 6139 17836 6184 17864
rect 2133 17799 2191 17805
rect 2133 17765 2145 17799
rect 2179 17796 2191 17799
rect 2746 17796 2774 17836
rect 3786 17796 3792 17808
rect 2179 17768 2774 17796
rect 3747 17768 3792 17796
rect 2179 17765 2191 17768
rect 2133 17759 2191 17765
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 5736 17796 5764 17836
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 8938 17864 8944 17876
rect 8899 17836 8944 17864
rect 8938 17824 8944 17836
rect 8996 17824 9002 17876
rect 13265 17867 13323 17873
rect 9048 17836 13124 17864
rect 9048 17796 9076 17836
rect 12618 17796 12624 17808
rect 5736 17768 9076 17796
rect 9140 17768 12624 17796
rect 9140 17728 9168 17768
rect 12618 17756 12624 17768
rect 12676 17756 12682 17808
rect 6840 17700 9168 17728
rect 1854 17660 1860 17672
rect 1815 17632 1860 17660
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 2682 17660 2688 17672
rect 2643 17632 2688 17660
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3384 17632 3985 17660
rect 3384 17620 3390 17632
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 3973 17623 4031 17629
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 6840 17669 6868 17700
rect 9490 17688 9496 17740
rect 9548 17688 9554 17740
rect 13096 17728 13124 17836
rect 13265 17833 13277 17867
rect 13311 17864 13323 17867
rect 13311 17836 15608 17864
rect 13311 17833 13323 17836
rect 13265 17827 13323 17833
rect 15580 17796 15608 17836
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15933 17867 15991 17873
rect 15933 17864 15945 17867
rect 15712 17836 15945 17864
rect 15712 17824 15718 17836
rect 15933 17833 15945 17836
rect 15979 17833 15991 17867
rect 15933 17827 15991 17833
rect 16206 17824 16212 17876
rect 16264 17864 16270 17876
rect 18141 17867 18199 17873
rect 18141 17864 18153 17867
rect 16264 17836 18153 17864
rect 16264 17824 16270 17836
rect 18141 17833 18153 17836
rect 18187 17833 18199 17867
rect 18141 17827 18199 17833
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 26234 17864 26240 17876
rect 18288 17836 26240 17864
rect 18288 17824 18294 17836
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 27154 17864 27160 17876
rect 27115 17836 27160 17864
rect 27154 17824 27160 17836
rect 27212 17824 27218 17876
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 29549 17867 29607 17873
rect 29549 17864 29561 17867
rect 29052 17836 29561 17864
rect 29052 17824 29058 17836
rect 29549 17833 29561 17836
rect 29595 17833 29607 17867
rect 29549 17827 29607 17833
rect 30282 17824 30288 17876
rect 30340 17864 30346 17876
rect 31478 17864 31484 17876
rect 30340 17836 31484 17864
rect 30340 17824 30346 17836
rect 31478 17824 31484 17836
rect 31536 17824 31542 17876
rect 37458 17864 37464 17876
rect 37200 17836 37464 17864
rect 21542 17796 21548 17808
rect 15580 17768 21548 17796
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 29917 17799 29975 17805
rect 29917 17796 29929 17799
rect 27264 17768 29929 17796
rect 18506 17728 18512 17740
rect 13096 17700 14679 17728
rect 18467 17700 18512 17728
rect 9385 17673 9443 17679
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 9122 17660 9128 17672
rect 9083 17632 9128 17660
rect 7101 17623 7159 17629
rect 5068 17595 5126 17601
rect 5068 17561 5080 17595
rect 5114 17592 5126 17595
rect 6641 17595 6699 17601
rect 6641 17592 6653 17595
rect 5114 17564 6653 17592
rect 5114 17561 5126 17564
rect 5068 17555 5126 17561
rect 6641 17561 6653 17564
rect 6687 17561 6699 17595
rect 6641 17555 6699 17561
rect 6730 17552 6736 17604
rect 6788 17592 6794 17604
rect 7116 17592 7144 17623
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9214 17620 9220 17672
rect 9272 17670 9278 17672
rect 9385 17670 9397 17673
rect 9272 17642 9397 17670
rect 9272 17620 9278 17642
rect 9385 17639 9397 17642
rect 9431 17639 9443 17673
rect 9385 17633 9443 17639
rect 9508 17656 9536 17688
rect 9674 17660 9680 17672
rect 9646 17656 9680 17660
rect 9508 17628 9680 17656
rect 9674 17620 9680 17628
rect 9732 17620 9738 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12250 17660 12256 17672
rect 12207 17632 12256 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12768 17632 12817 17660
rect 12768 17620 12774 17632
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 13354 17660 13360 17672
rect 13127 17632 13360 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 13872 17632 14565 17660
rect 13872 17620 13878 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14651 17660 14679 17700
rect 18506 17688 18512 17700
rect 18564 17688 18570 17740
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18840 17700 19257 17728
rect 18840 17688 18846 17700
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 23934 17688 23940 17740
rect 23992 17728 23998 17740
rect 24394 17728 24400 17740
rect 23992 17700 24400 17728
rect 23992 17688 23998 17700
rect 24394 17688 24400 17700
rect 24452 17688 24458 17740
rect 27264 17737 27292 17768
rect 29917 17765 29929 17768
rect 29963 17765 29975 17799
rect 29917 17759 29975 17765
rect 32030 17756 32036 17808
rect 32088 17756 32094 17808
rect 27249 17731 27307 17737
rect 27249 17697 27261 17731
rect 27295 17697 27307 17731
rect 27249 17691 27307 17697
rect 27430 17688 27436 17740
rect 27488 17728 27494 17740
rect 31202 17728 31208 17740
rect 27488 17700 31208 17728
rect 27488 17688 27494 17700
rect 31202 17688 31208 17700
rect 31260 17728 31266 17740
rect 31846 17728 31852 17740
rect 31260 17700 31852 17728
rect 31260 17688 31266 17700
rect 31846 17688 31852 17700
rect 31904 17688 31910 17740
rect 32048 17728 32076 17756
rect 32309 17731 32367 17737
rect 32309 17728 32321 17731
rect 32048 17700 32321 17728
rect 32309 17697 32321 17700
rect 32355 17697 32367 17731
rect 32309 17691 32367 17697
rect 16114 17660 16120 17672
rect 14651 17632 16120 17660
rect 14553 17623 14611 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 18322 17660 18328 17672
rect 18283 17632 18328 17660
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18414 17620 18420 17672
rect 18472 17660 18478 17672
rect 18601 17663 18659 17669
rect 18472 17632 18517 17660
rect 18472 17620 18478 17632
rect 18601 17629 18613 17663
rect 18647 17660 18659 17663
rect 18690 17660 18696 17672
rect 18647 17632 18696 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 19978 17660 19984 17672
rect 19567 17632 19984 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 21634 17660 21640 17672
rect 21595 17632 21640 17660
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 26973 17663 27031 17669
rect 26973 17629 26985 17663
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 6788 17564 7144 17592
rect 6788 17552 6794 17564
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 12986 17592 12992 17604
rect 9364 17564 9409 17592
rect 9646 17564 12434 17592
rect 12947 17564 12992 17592
rect 9364 17552 9370 17564
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 7009 17527 7067 17533
rect 7009 17524 7021 17527
rect 6236 17496 7021 17524
rect 6236 17484 6242 17496
rect 7009 17493 7021 17496
rect 7055 17493 7067 17527
rect 7009 17487 7067 17493
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 9122 17524 9128 17536
rect 7524 17496 9128 17524
rect 7524 17484 7530 17496
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 9490 17484 9496 17536
rect 9548 17524 9554 17536
rect 9646 17524 9674 17564
rect 9548 17496 9674 17524
rect 9548 17484 9554 17496
rect 12158 17484 12164 17536
rect 12216 17524 12222 17536
rect 12253 17527 12311 17533
rect 12253 17524 12265 17527
rect 12216 17496 12265 17524
rect 12216 17484 12222 17496
rect 12253 17493 12265 17496
rect 12299 17493 12311 17527
rect 12406 17524 12434 17564
rect 12986 17552 12992 17564
rect 13044 17552 13050 17604
rect 14820 17595 14878 17601
rect 14820 17561 14832 17595
rect 14866 17592 14878 17595
rect 15286 17592 15292 17604
rect 14866 17564 15292 17592
rect 14866 17561 14878 17564
rect 14820 17555 14878 17561
rect 15286 17552 15292 17564
rect 15344 17552 15350 17604
rect 17126 17552 17132 17604
rect 17184 17592 17190 17604
rect 21910 17601 21916 17604
rect 17184 17564 18276 17592
rect 17184 17552 17190 17564
rect 14734 17524 14740 17536
rect 12406 17496 14740 17524
rect 12253 17487 12311 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 18138 17524 18144 17536
rect 15160 17496 18144 17524
rect 15160 17484 15166 17496
rect 18138 17484 18144 17496
rect 18196 17484 18202 17536
rect 18248 17524 18276 17564
rect 21904 17555 21916 17601
rect 21968 17592 21974 17604
rect 24670 17601 24676 17604
rect 21968 17564 22004 17592
rect 21910 17552 21916 17555
rect 21968 17552 21974 17564
rect 24664 17555 24676 17601
rect 24728 17592 24734 17604
rect 26988 17592 27016 17623
rect 27062 17620 27068 17672
rect 27120 17660 27126 17672
rect 29546 17660 29552 17672
rect 27120 17632 27165 17660
rect 29507 17632 29552 17660
rect 27120 17620 27126 17632
rect 29546 17620 29552 17632
rect 29604 17620 29610 17672
rect 29733 17663 29791 17669
rect 29733 17629 29745 17663
rect 29779 17660 29791 17663
rect 30558 17660 30564 17672
rect 29779 17632 30564 17660
rect 29779 17629 29791 17632
rect 29733 17623 29791 17629
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 32033 17663 32091 17669
rect 32033 17629 32045 17663
rect 32079 17660 32091 17663
rect 32398 17660 32404 17672
rect 32079 17632 32404 17660
rect 32079 17629 32091 17632
rect 32033 17623 32091 17629
rect 32398 17620 32404 17632
rect 32456 17660 32462 17672
rect 34701 17663 34759 17669
rect 34701 17660 34713 17663
rect 32456 17632 34713 17660
rect 32456 17620 32462 17632
rect 34701 17629 34713 17632
rect 34747 17660 34759 17663
rect 34790 17660 34796 17672
rect 34747 17632 34796 17660
rect 34747 17629 34759 17632
rect 34701 17623 34759 17629
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 37200 17669 37228 17836
rect 37458 17824 37464 17836
rect 37516 17824 37522 17876
rect 39853 17867 39911 17873
rect 39853 17833 39865 17867
rect 39899 17864 39911 17867
rect 40034 17864 40040 17876
rect 39899 17836 40040 17864
rect 39899 17833 39911 17836
rect 39853 17827 39911 17833
rect 40034 17824 40040 17836
rect 40092 17824 40098 17876
rect 48314 17864 48320 17876
rect 42628 17836 45508 17864
rect 48275 17836 48320 17864
rect 38010 17728 38016 17740
rect 37292 17700 38016 17728
rect 37292 17669 37320 17700
rect 38010 17688 38016 17700
rect 38068 17688 38074 17740
rect 40494 17688 40500 17740
rect 40552 17728 40558 17740
rect 41046 17728 41052 17740
rect 40552 17700 41052 17728
rect 40552 17688 40558 17700
rect 41046 17688 41052 17700
rect 41104 17728 41110 17740
rect 42628 17737 42656 17836
rect 45480 17737 45508 17836
rect 48314 17824 48320 17836
rect 48372 17864 48378 17876
rect 48590 17864 48596 17876
rect 48372 17836 48596 17864
rect 48372 17824 48378 17836
rect 48590 17824 48596 17836
rect 48648 17824 48654 17876
rect 42613 17731 42671 17737
rect 42613 17728 42625 17731
rect 41104 17700 42625 17728
rect 41104 17688 41110 17700
rect 42613 17697 42625 17700
rect 42659 17697 42671 17731
rect 42613 17691 42671 17697
rect 45465 17731 45523 17737
rect 45465 17697 45477 17731
rect 45511 17697 45523 17731
rect 45465 17691 45523 17697
rect 37185 17663 37243 17669
rect 37185 17629 37197 17663
rect 37231 17629 37243 17663
rect 37185 17623 37243 17629
rect 37277 17663 37335 17669
rect 37277 17629 37289 17663
rect 37323 17629 37335 17663
rect 37277 17623 37335 17629
rect 37366 17620 37372 17672
rect 37424 17660 37430 17672
rect 37553 17663 37611 17669
rect 37424 17632 37469 17660
rect 37424 17620 37430 17632
rect 37553 17629 37565 17663
rect 37599 17629 37611 17663
rect 40034 17660 40040 17672
rect 39995 17632 40040 17660
rect 37553 17623 37611 17629
rect 33686 17592 33692 17604
rect 24728 17564 24764 17592
rect 26988 17564 33692 17592
rect 24670 17552 24676 17555
rect 24728 17552 24734 17564
rect 33686 17552 33692 17564
rect 33744 17552 33750 17604
rect 34054 17552 34060 17604
rect 34112 17592 34118 17604
rect 37568 17592 37596 17623
rect 40034 17620 40040 17632
rect 40092 17620 40098 17672
rect 40310 17660 40316 17672
rect 40271 17632 40316 17660
rect 40310 17620 40316 17632
rect 40368 17620 40374 17672
rect 41386 17632 44128 17660
rect 41386 17592 41414 17632
rect 42886 17601 42892 17604
rect 34112 17564 41414 17592
rect 34112 17552 34118 17564
rect 42880 17555 42892 17601
rect 42944 17592 42950 17604
rect 42944 17564 42980 17592
rect 42886 17552 42892 17555
rect 42944 17552 42950 17564
rect 20622 17524 20628 17536
rect 18248 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 22370 17484 22376 17536
rect 22428 17524 22434 17536
rect 23017 17527 23075 17533
rect 23017 17524 23029 17527
rect 22428 17496 23029 17524
rect 22428 17484 22434 17496
rect 23017 17493 23029 17496
rect 23063 17493 23075 17527
rect 23017 17487 23075 17493
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 25280 17496 25789 17524
rect 25280 17484 25286 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 25777 17487 25835 17493
rect 34698 17484 34704 17536
rect 34756 17524 34762 17536
rect 34885 17527 34943 17533
rect 34885 17524 34897 17527
rect 34756 17496 34897 17524
rect 34756 17484 34762 17496
rect 34885 17493 34897 17496
rect 34931 17524 34943 17527
rect 35986 17524 35992 17536
rect 34931 17496 35992 17524
rect 34931 17493 34943 17496
rect 34885 17487 34943 17493
rect 35986 17484 35992 17496
rect 36044 17484 36050 17536
rect 36909 17527 36967 17533
rect 36909 17493 36921 17527
rect 36955 17524 36967 17527
rect 37182 17524 37188 17536
rect 36955 17496 37188 17524
rect 36955 17493 36967 17496
rect 36909 17487 36967 17493
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 39850 17484 39856 17536
rect 39908 17524 39914 17536
rect 40221 17527 40279 17533
rect 40221 17524 40233 17527
rect 39908 17496 40233 17524
rect 39908 17484 39914 17496
rect 40221 17493 40233 17496
rect 40267 17493 40279 17527
rect 43990 17524 43996 17536
rect 43951 17496 43996 17524
rect 40221 17487 40279 17493
rect 43990 17484 43996 17496
rect 44048 17484 44054 17536
rect 44100 17524 44128 17632
rect 45278 17552 45284 17604
rect 45336 17592 45342 17604
rect 45710 17595 45768 17601
rect 45710 17592 45722 17595
rect 45336 17564 45722 17592
rect 45336 17552 45342 17564
rect 45710 17561 45722 17564
rect 45756 17561 45768 17595
rect 47854 17592 47860 17604
rect 45710 17555 45768 17561
rect 46768 17564 47860 17592
rect 46768 17524 46796 17564
rect 47854 17552 47860 17564
rect 47912 17592 47918 17604
rect 48225 17595 48283 17601
rect 48225 17592 48237 17595
rect 47912 17564 48237 17592
rect 47912 17552 47918 17564
rect 48225 17561 48237 17564
rect 48271 17561 48283 17595
rect 48225 17555 48283 17561
rect 44100 17496 46796 17524
rect 46845 17527 46903 17533
rect 46845 17493 46857 17527
rect 46891 17524 46903 17527
rect 47118 17524 47124 17536
rect 46891 17496 47124 17524
rect 46891 17493 46903 17496
rect 46845 17487 46903 17493
rect 47118 17484 47124 17496
rect 47176 17484 47182 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 15102 17320 15108 17332
rect 6880 17292 15108 17320
rect 6880 17280 6886 17292
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 15286 17320 15292 17332
rect 15247 17292 15292 17320
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15654 17320 15660 17332
rect 15615 17292 15660 17320
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 22186 17320 22192 17332
rect 16172 17292 22192 17320
rect 16172 17280 16178 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22370 17320 22376 17332
rect 22331 17292 22376 17320
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 24670 17320 24676 17332
rect 24631 17292 24676 17320
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 25498 17320 25504 17332
rect 24780 17292 25504 17320
rect 1946 17212 1952 17264
rect 2004 17252 2010 17264
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 2004 17224 3464 17252
rect 2004 17212 2010 17224
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1412 17116 1440 17147
rect 2406 17144 2412 17196
rect 2464 17184 2470 17196
rect 2685 17187 2743 17193
rect 2685 17184 2697 17187
rect 2464 17156 2697 17184
rect 2464 17144 2470 17156
rect 2685 17153 2697 17156
rect 2731 17153 2743 17187
rect 3326 17184 3332 17196
rect 3287 17156 3332 17184
rect 2685 17147 2743 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 3436 17184 3464 17224
rect 6840 17224 13277 17252
rect 6840 17184 6868 17224
rect 13265 17221 13277 17224
rect 13311 17221 13323 17255
rect 13265 17215 13323 17221
rect 13817 17255 13875 17261
rect 13817 17221 13829 17255
rect 13863 17252 13875 17255
rect 13863 17224 15424 17252
rect 13863 17221 13875 17224
rect 13817 17215 13875 17221
rect 15396 17196 15424 17224
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 24780 17252 24808 17292
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 26237 17323 26295 17329
rect 26237 17289 26249 17323
rect 26283 17320 26295 17323
rect 27062 17320 27068 17332
rect 26283 17292 27068 17320
rect 26283 17289 26295 17292
rect 26237 17283 26295 17289
rect 26252 17252 26280 17283
rect 27062 17280 27068 17292
rect 27120 17280 27126 17332
rect 30282 17280 30288 17332
rect 30340 17320 30346 17332
rect 31573 17323 31631 17329
rect 31573 17320 31585 17323
rect 30340 17292 31585 17320
rect 30340 17280 30346 17292
rect 31573 17289 31585 17292
rect 31619 17289 31631 17323
rect 31573 17283 31631 17289
rect 32674 17280 32680 17332
rect 32732 17280 32738 17332
rect 38930 17320 38936 17332
rect 38891 17292 38936 17320
rect 38930 17280 38936 17292
rect 38988 17280 38994 17332
rect 42886 17320 42892 17332
rect 42847 17292 42892 17320
rect 42886 17280 42892 17292
rect 42944 17280 42950 17332
rect 45278 17320 45284 17332
rect 45239 17292 45284 17320
rect 45278 17280 45284 17292
rect 45336 17280 45342 17332
rect 18472 17224 24808 17252
rect 25148 17224 26280 17252
rect 27617 17255 27675 17261
rect 18472 17212 18478 17224
rect 3436 17156 6868 17184
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 7834 17184 7840 17196
rect 7791 17156 7840 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8012 17187 8070 17193
rect 8012 17153 8024 17187
rect 8058 17184 8070 17187
rect 8938 17184 8944 17196
rect 8058 17156 8944 17184
rect 8058 17153 8070 17156
rect 8012 17147 8070 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 10134 17184 10140 17196
rect 9180 17156 10140 17184
rect 9180 17144 9186 17156
rect 10134 17144 10140 17156
rect 10192 17144 10198 17196
rect 12158 17184 12164 17196
rect 12119 17156 12164 17184
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 12342 17184 12348 17196
rect 12303 17156 12348 17184
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 13354 17184 13360 17196
rect 13315 17156 13360 17184
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 6638 17116 6644 17128
rect 1412 17088 6644 17116
rect 6638 17076 6644 17088
rect 6696 17076 6702 17128
rect 14384 17116 14412 17147
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 15436 17156 15485 17184
rect 15436 17144 15442 17156
rect 15473 17153 15485 17156
rect 15519 17153 15531 17187
rect 15473 17147 15531 17153
rect 15749 17187 15807 17193
rect 15749 17153 15761 17187
rect 15795 17184 15807 17187
rect 18506 17184 18512 17196
rect 15795 17156 18512 17184
rect 15795 17153 15807 17156
rect 15749 17147 15807 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17184 19027 17187
rect 19058 17184 19064 17196
rect 19015 17156 19064 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 22189 17187 22247 17193
rect 22189 17184 22201 17187
rect 19208 17156 22201 17184
rect 19208 17144 19214 17156
rect 22189 17153 22201 17156
rect 22235 17184 22247 17187
rect 22278 17184 22284 17196
rect 22235 17156 22284 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22646 17184 22652 17196
rect 22511 17156 22652 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 24949 17190 25007 17193
rect 25148 17190 25176 17224
rect 27617 17221 27629 17255
rect 27663 17252 27675 17255
rect 28902 17252 28908 17264
rect 27663 17224 28908 17252
rect 27663 17221 27675 17224
rect 27617 17215 27675 17221
rect 28902 17212 28908 17224
rect 28960 17252 28966 17264
rect 31205 17255 31263 17261
rect 31205 17252 31217 17255
rect 28960 17224 31217 17252
rect 28960 17212 28966 17224
rect 31205 17221 31217 17224
rect 31251 17221 31263 17255
rect 31205 17215 31263 17221
rect 31846 17212 31852 17264
rect 31904 17252 31910 17264
rect 32401 17255 32459 17261
rect 32401 17252 32413 17255
rect 31904 17224 32413 17252
rect 31904 17212 31910 17224
rect 32401 17221 32413 17224
rect 32447 17221 32459 17255
rect 32401 17215 32459 17221
rect 32493 17255 32551 17261
rect 32493 17221 32505 17255
rect 32539 17252 32551 17255
rect 32692 17252 32720 17280
rect 32539 17224 32720 17252
rect 32539 17221 32551 17224
rect 32493 17215 32551 17221
rect 24949 17187 25176 17190
rect 24949 17153 24961 17187
rect 24995 17162 25176 17187
rect 26050 17184 26056 17196
rect 24995 17153 25007 17162
rect 26011 17156 26056 17184
rect 24949 17147 25007 17153
rect 26050 17144 26056 17156
rect 26108 17144 26114 17196
rect 26234 17144 26240 17196
rect 26292 17184 26298 17196
rect 26878 17184 26884 17196
rect 26292 17156 26884 17184
rect 26292 17144 26298 17156
rect 26878 17144 26884 17156
rect 26936 17144 26942 17196
rect 27430 17184 27436 17196
rect 27391 17156 27436 17184
rect 27430 17144 27436 17156
rect 27488 17144 27494 17196
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 29822 17184 29828 17196
rect 27580 17156 29828 17184
rect 27580 17144 27586 17156
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 30926 17184 30932 17196
rect 30887 17156 30932 17184
rect 30926 17144 30932 17156
rect 30984 17144 30990 17196
rect 31110 17193 31116 17196
rect 31077 17187 31116 17193
rect 31077 17153 31089 17187
rect 31077 17147 31116 17153
rect 31110 17144 31116 17147
rect 31168 17144 31174 17196
rect 31294 17184 31300 17196
rect 31255 17156 31300 17184
rect 31294 17144 31300 17156
rect 31352 17144 31358 17196
rect 31394 17187 31452 17193
rect 31394 17153 31406 17187
rect 31440 17184 31452 17187
rect 31440 17156 31524 17184
rect 31440 17153 31452 17156
rect 31394 17147 31452 17153
rect 12268 17088 14412 17116
rect 12268 17060 12296 17088
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 17184 17088 17417 17116
rect 17184 17076 17190 17088
rect 17405 17085 17417 17088
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 17681 17119 17739 17125
rect 17681 17116 17693 17119
rect 17552 17088 17693 17116
rect 17552 17076 17558 17088
rect 17681 17085 17693 17088
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 18598 17076 18604 17128
rect 18656 17116 18662 17128
rect 18693 17119 18751 17125
rect 18693 17116 18705 17119
rect 18656 17088 18705 17116
rect 18656 17076 18662 17088
rect 18693 17085 18705 17088
rect 18739 17085 18751 17119
rect 18693 17079 18751 17085
rect 21910 17076 21916 17128
rect 21968 17116 21974 17128
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21968 17088 22017 17116
rect 21968 17076 21974 17088
rect 22005 17085 22017 17088
rect 22051 17085 22063 17119
rect 22005 17079 22063 17085
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 24857 17119 24915 17125
rect 22152 17088 24808 17116
rect 22152 17076 22158 17088
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 11974 17048 11980 17060
rect 1728 17020 7604 17048
rect 1728 17008 1734 17020
rect 1394 16940 1400 16992
rect 1452 16980 1458 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 1452 16952 1593 16980
rect 1452 16940 1458 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 2498 16980 2504 16992
rect 2459 16952 2504 16980
rect 1581 16943 1639 16949
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 3145 16983 3203 16989
rect 3145 16949 3157 16983
rect 3191 16980 3203 16983
rect 7466 16980 7472 16992
rect 3191 16952 7472 16980
rect 3191 16949 3203 16952
rect 3145 16943 3203 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 7576 16980 7604 17020
rect 8680 17020 11980 17048
rect 8680 16980 8708 17020
rect 11974 17008 11980 17020
rect 12032 17008 12038 17060
rect 12250 17008 12256 17060
rect 12308 17008 12314 17060
rect 12345 17051 12403 17057
rect 12345 17017 12357 17051
rect 12391 17048 12403 17051
rect 24670 17048 24676 17060
rect 12391 17020 24676 17048
rect 12391 17017 12403 17020
rect 12345 17011 12403 17017
rect 24670 17008 24676 17020
rect 24728 17008 24734 17060
rect 24780 17048 24808 17088
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 25038 17116 25044 17128
rect 24903 17088 25044 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 25038 17076 25044 17088
rect 25096 17076 25102 17128
rect 25222 17116 25228 17128
rect 25135 17088 25228 17116
rect 25222 17076 25228 17088
rect 25280 17076 25286 17128
rect 25314 17076 25320 17128
rect 25372 17116 25378 17128
rect 25372 17088 25417 17116
rect 25372 17076 25378 17088
rect 25498 17076 25504 17128
rect 25556 17116 25562 17128
rect 30282 17116 30288 17128
rect 25556 17088 30288 17116
rect 25556 17076 25562 17088
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 31496 17116 31524 17156
rect 32030 17144 32036 17196
rect 32088 17184 32094 17196
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 32088 17156 32137 17184
rect 32088 17144 32094 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32214 17144 32220 17196
rect 32272 17184 32278 17196
rect 32631 17187 32689 17193
rect 32272 17156 32317 17184
rect 32272 17144 32278 17156
rect 32631 17153 32643 17187
rect 32677 17184 32689 17187
rect 32766 17184 32772 17196
rect 32677 17156 32772 17184
rect 32677 17153 32689 17156
rect 32631 17147 32689 17153
rect 31662 17116 31668 17128
rect 31496 17088 31668 17116
rect 31662 17076 31668 17088
rect 31720 17116 31726 17128
rect 32646 17116 32674 17147
rect 32766 17144 32772 17156
rect 32824 17144 32830 17196
rect 37274 17144 37280 17196
rect 37332 17184 37338 17196
rect 37809 17187 37867 17193
rect 37809 17184 37821 17187
rect 37332 17156 37821 17184
rect 37332 17144 37338 17156
rect 37809 17153 37821 17156
rect 37855 17153 37867 17187
rect 43070 17184 43076 17196
rect 43031 17156 43076 17184
rect 37809 17147 37867 17153
rect 43070 17144 43076 17156
rect 43128 17144 43134 17196
rect 45465 17187 45523 17193
rect 45465 17153 45477 17187
rect 45511 17184 45523 17187
rect 45554 17184 45560 17196
rect 45511 17156 45560 17184
rect 45511 17153 45523 17156
rect 45465 17147 45523 17153
rect 45554 17144 45560 17156
rect 45612 17144 45618 17196
rect 31720 17088 32674 17116
rect 31720 17076 31726 17088
rect 37366 17076 37372 17128
rect 37424 17116 37430 17128
rect 37553 17119 37611 17125
rect 37553 17116 37565 17119
rect 37424 17088 37565 17116
rect 37424 17076 37430 17088
rect 37553 17085 37565 17088
rect 37599 17085 37611 17119
rect 37553 17079 37611 17085
rect 25240 17048 25268 17076
rect 24780 17020 25268 17048
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 32769 17051 32827 17057
rect 32769 17048 32781 17051
rect 25740 17020 32781 17048
rect 25740 17008 25746 17020
rect 32769 17017 32781 17020
rect 32815 17017 32827 17051
rect 32769 17011 32827 17017
rect 9122 16980 9128 16992
rect 7576 16952 8708 16980
rect 9083 16952 9128 16980
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12768 16952 13093 16980
rect 12768 16940 12774 16952
rect 13081 16949 13093 16952
rect 13127 16980 13139 16983
rect 13906 16980 13912 16992
rect 13127 16952 13912 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14458 16980 14464 16992
rect 14419 16952 14464 16980
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 40034 16980 40040 16992
rect 15436 16952 40040 16980
rect 15436 16940 15442 16952
rect 40034 16940 40040 16952
rect 40092 16940 40098 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 8938 16776 8944 16788
rect 2096 16748 7604 16776
rect 8899 16748 8944 16776
rect 2096 16736 2102 16748
rect 7576 16708 7604 16748
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 12250 16776 12256 16788
rect 9048 16748 11933 16776
rect 12211 16748 12256 16776
rect 9048 16708 9076 16748
rect 7576 16680 9076 16708
rect 9214 16640 9220 16652
rect 8312 16612 9220 16640
rect 1486 16532 1492 16584
rect 1544 16572 1550 16584
rect 1857 16575 1915 16581
rect 1857 16572 1869 16575
rect 1544 16544 1869 16572
rect 1544 16532 1550 16544
rect 1857 16541 1869 16544
rect 1903 16572 1915 16575
rect 1946 16572 1952 16584
rect 1903 16544 1952 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2124 16575 2182 16581
rect 2124 16541 2136 16575
rect 2170 16572 2182 16575
rect 2498 16572 2504 16584
rect 2170 16544 2504 16572
rect 2170 16541 2182 16544
rect 2124 16535 2182 16541
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 3970 16572 3976 16584
rect 3931 16544 3976 16572
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 4890 16504 4896 16516
rect 3252 16476 4896 16504
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 3252 16445 3280 16476
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 8110 16464 8116 16516
rect 8168 16504 8174 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 8168 16476 8217 16504
rect 8168 16464 8174 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 3237 16439 3295 16445
rect 3237 16436 3249 16439
rect 2832 16408 3249 16436
rect 2832 16396 2838 16408
rect 3237 16405 3249 16408
rect 3283 16405 3295 16439
rect 3786 16436 3792 16448
rect 3747 16408 3792 16436
rect 3237 16399 3295 16405
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 6730 16396 6736 16448
rect 6788 16436 6794 16448
rect 8312 16445 8340 16612
rect 9214 16600 9220 16612
rect 9272 16640 9278 16652
rect 10870 16640 10876 16652
rect 9272 16612 9444 16640
rect 10831 16612 10876 16640
rect 9272 16600 9278 16612
rect 9416 16581 9444 16612
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 11905 16640 11933 16748
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 14642 16776 14648 16788
rect 14603 16748 14648 16776
rect 14642 16736 14648 16748
rect 14700 16736 14706 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 17034 16776 17040 16788
rect 14792 16748 17040 16776
rect 14792 16736 14798 16748
rect 17034 16736 17040 16748
rect 17092 16736 17098 16788
rect 35253 16779 35311 16785
rect 35253 16776 35265 16779
rect 17236 16748 35265 16776
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 12986 16708 12992 16720
rect 12032 16680 12992 16708
rect 12032 16668 12038 16680
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 13354 16708 13360 16720
rect 13315 16680 13360 16708
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 17236 16640 17264 16748
rect 35253 16745 35265 16748
rect 35299 16776 35311 16779
rect 35618 16776 35624 16788
rect 35299 16748 35624 16776
rect 35299 16745 35311 16748
rect 35253 16739 35311 16745
rect 35618 16736 35624 16748
rect 35676 16776 35682 16788
rect 35805 16779 35863 16785
rect 35805 16776 35817 16779
rect 35676 16748 35817 16776
rect 35676 16736 35682 16748
rect 35805 16745 35817 16748
rect 35851 16745 35863 16779
rect 35805 16739 35863 16745
rect 42889 16779 42947 16785
rect 42889 16745 42901 16779
rect 42935 16745 42947 16779
rect 43070 16776 43076 16788
rect 43031 16748 43076 16776
rect 42889 16739 42947 16745
rect 18874 16668 18880 16720
rect 18932 16708 18938 16720
rect 22094 16708 22100 16720
rect 18932 16680 22100 16708
rect 18932 16668 18938 16680
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 24670 16668 24676 16720
rect 24728 16708 24734 16720
rect 27430 16708 27436 16720
rect 24728 16680 27436 16708
rect 24728 16668 24734 16680
rect 27430 16668 27436 16680
rect 27488 16668 27494 16720
rect 29362 16668 29368 16720
rect 29420 16708 29426 16720
rect 31846 16708 31852 16720
rect 29420 16680 31852 16708
rect 29420 16668 29426 16680
rect 31846 16668 31852 16680
rect 31904 16668 31910 16720
rect 32858 16668 32864 16720
rect 32916 16708 32922 16720
rect 42904 16708 42932 16739
rect 43070 16736 43076 16748
rect 43128 16736 43134 16788
rect 45554 16736 45560 16788
rect 45612 16776 45618 16788
rect 45612 16748 45657 16776
rect 45612 16736 45618 16748
rect 32916 16680 37320 16708
rect 32916 16668 32922 16680
rect 11905 16612 17264 16640
rect 18417 16643 18475 16649
rect 18417 16609 18429 16643
rect 18463 16640 18475 16643
rect 18463 16612 19334 16640
rect 18463 16609 18475 16612
rect 18417 16603 18475 16609
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16541 9459 16575
rect 18322 16572 18328 16584
rect 18283 16544 18328 16572
rect 9401 16535 9459 16541
rect 9140 16504 9168 16535
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 18432 16544 18521 16572
rect 18432 16516 18460 16544
rect 18509 16541 18521 16544
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16572 18659 16575
rect 18690 16572 18696 16584
rect 18647 16544 18696 16572
rect 18647 16541 18659 16544
rect 18601 16535 18659 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19306 16572 19334 16612
rect 22186 16600 22192 16652
rect 22244 16640 22250 16652
rect 22244 16612 24532 16640
rect 22244 16600 22250 16612
rect 24118 16572 24124 16584
rect 19306 16544 24124 16572
rect 24118 16532 24124 16544
rect 24176 16532 24182 16584
rect 24504 16572 24532 16612
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 36909 16643 36967 16649
rect 36909 16640 36921 16643
rect 26108 16612 36921 16640
rect 26108 16600 26114 16612
rect 36909 16609 36921 16612
rect 36955 16609 36967 16643
rect 36909 16603 36967 16609
rect 36998 16600 37004 16652
rect 37056 16640 37062 16652
rect 37182 16640 37188 16652
rect 37056 16612 37101 16640
rect 37143 16612 37188 16640
rect 37056 16600 37062 16612
rect 37182 16600 37188 16612
rect 37240 16600 37246 16652
rect 24854 16572 24860 16584
rect 24504 16544 24860 16572
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 25130 16572 25136 16584
rect 25043 16544 25136 16572
rect 25130 16532 25136 16544
rect 25188 16572 25194 16584
rect 26142 16572 26148 16584
rect 25188 16544 26148 16572
rect 25188 16532 25194 16544
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 26568 16544 29960 16572
rect 26568 16532 26574 16544
rect 9140 16476 9444 16504
rect 8297 16439 8355 16445
rect 8297 16436 8309 16439
rect 6788 16408 8309 16436
rect 6788 16396 6794 16408
rect 8297 16405 8309 16408
rect 8343 16405 8355 16439
rect 8297 16399 8355 16405
rect 9122 16396 9128 16448
rect 9180 16436 9186 16448
rect 9309 16439 9367 16445
rect 9309 16436 9321 16439
rect 9180 16408 9321 16436
rect 9180 16396 9186 16408
rect 9309 16405 9321 16408
rect 9355 16405 9367 16439
rect 9416 16436 9444 16476
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 11118 16507 11176 16513
rect 11118 16504 11130 16507
rect 10836 16476 11130 16504
rect 10836 16464 10842 16476
rect 11118 16473 11130 16476
rect 11164 16473 11176 16507
rect 11118 16467 11176 16473
rect 13078 16464 13084 16516
rect 13136 16504 13142 16516
rect 13173 16507 13231 16513
rect 13173 16504 13185 16507
rect 13136 16476 13185 16504
rect 13136 16464 13142 16476
rect 13173 16473 13185 16476
rect 13219 16473 13231 16507
rect 14550 16504 14556 16516
rect 14511 16476 14556 16504
rect 13173 16467 13231 16473
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 15436 16476 18276 16504
rect 15436 16464 15442 16476
rect 10870 16436 10876 16448
rect 9416 16408 10876 16436
rect 9309 16399 9367 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 18141 16439 18199 16445
rect 18141 16436 18153 16439
rect 12676 16408 18153 16436
rect 12676 16396 12682 16408
rect 18141 16405 18153 16408
rect 18187 16405 18199 16439
rect 18248 16436 18276 16476
rect 18414 16464 18420 16516
rect 18472 16464 18478 16516
rect 29362 16504 29368 16516
rect 18524 16476 29368 16504
rect 18524 16436 18552 16476
rect 29362 16464 29368 16476
rect 29420 16464 29426 16516
rect 29546 16504 29552 16516
rect 29507 16476 29552 16504
rect 29546 16464 29552 16476
rect 29604 16464 29610 16516
rect 29733 16507 29791 16513
rect 29733 16473 29745 16507
rect 29779 16504 29791 16507
rect 29822 16504 29828 16516
rect 29779 16476 29828 16504
rect 29779 16473 29791 16476
rect 29733 16467 29791 16473
rect 29822 16464 29828 16476
rect 29880 16464 29886 16516
rect 29932 16504 29960 16544
rect 30374 16532 30380 16584
rect 30432 16572 30438 16584
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 30432 16544 30757 16572
rect 30432 16532 30438 16544
rect 30745 16541 30757 16544
rect 30791 16541 30803 16575
rect 30926 16572 30932 16584
rect 30887 16544 30932 16572
rect 30745 16535 30803 16541
rect 30926 16532 30932 16544
rect 30984 16532 30990 16584
rect 33778 16572 33784 16584
rect 33739 16544 33784 16572
rect 33778 16532 33784 16544
rect 33836 16532 33842 16584
rect 33962 16572 33968 16584
rect 33923 16544 33968 16572
rect 33962 16532 33968 16544
rect 34020 16532 34026 16584
rect 37093 16575 37151 16581
rect 35084 16544 36124 16572
rect 31202 16504 31208 16516
rect 29932 16476 31208 16504
rect 31202 16464 31208 16476
rect 31260 16464 31266 16516
rect 34790 16464 34796 16516
rect 34848 16504 34854 16516
rect 35084 16513 35112 16544
rect 35069 16507 35127 16513
rect 35069 16504 35081 16507
rect 34848 16476 35081 16504
rect 34848 16464 34854 16476
rect 35069 16473 35081 16476
rect 35115 16473 35127 16507
rect 35069 16467 35127 16473
rect 35253 16507 35311 16513
rect 35253 16473 35265 16507
rect 35299 16504 35311 16507
rect 35986 16504 35992 16516
rect 35299 16476 35992 16504
rect 35299 16473 35311 16476
rect 35253 16467 35311 16473
rect 35986 16464 35992 16476
rect 36044 16464 36050 16516
rect 36096 16504 36124 16544
rect 37093 16541 37105 16575
rect 37139 16572 37151 16575
rect 37292 16572 37320 16680
rect 42904 16680 44220 16708
rect 37366 16600 37372 16652
rect 37424 16640 37430 16652
rect 40218 16640 40224 16652
rect 37424 16612 40224 16640
rect 37424 16600 37430 16612
rect 40218 16600 40224 16612
rect 40276 16600 40282 16652
rect 40497 16643 40555 16649
rect 40497 16609 40509 16643
rect 40543 16640 40555 16643
rect 42904 16640 42932 16680
rect 40543 16612 42932 16640
rect 40543 16609 40555 16612
rect 40497 16603 40555 16609
rect 40512 16572 40540 16603
rect 43254 16600 43260 16652
rect 43312 16640 43318 16652
rect 43901 16643 43959 16649
rect 43901 16640 43913 16643
rect 43312 16612 43913 16640
rect 43312 16600 43318 16612
rect 43901 16609 43913 16612
rect 43947 16609 43959 16643
rect 43901 16603 43959 16609
rect 43990 16600 43996 16652
rect 44048 16640 44054 16652
rect 44048 16612 44093 16640
rect 44048 16600 44054 16612
rect 37139 16544 37320 16572
rect 37936 16544 40540 16572
rect 37139 16541 37151 16544
rect 37093 16535 37151 16541
rect 37936 16504 37964 16544
rect 40586 16532 40592 16584
rect 40644 16572 40650 16584
rect 41141 16575 41199 16581
rect 41141 16572 41153 16575
rect 40644 16544 41153 16572
rect 40644 16532 40650 16544
rect 41141 16541 41153 16544
rect 41187 16541 41199 16575
rect 43714 16572 43720 16584
rect 43675 16544 43720 16572
rect 41141 16535 41199 16541
rect 43714 16532 43720 16544
rect 43772 16532 43778 16584
rect 43806 16532 43812 16584
rect 43864 16572 43870 16584
rect 44192 16572 44220 16680
rect 45002 16640 45008 16652
rect 44963 16612 45008 16640
rect 45002 16600 45008 16612
rect 45060 16640 45066 16652
rect 45462 16640 45468 16652
rect 45060 16612 45468 16640
rect 45060 16600 45066 16612
rect 45462 16600 45468 16612
rect 45520 16600 45526 16652
rect 46400 16612 46704 16640
rect 45189 16575 45247 16581
rect 45189 16572 45201 16575
rect 43864 16544 43909 16572
rect 44192 16544 45201 16572
rect 43864 16532 43870 16544
rect 45189 16541 45201 16544
rect 45235 16572 45247 16575
rect 46400 16572 46428 16612
rect 46566 16572 46572 16584
rect 45235 16544 46428 16572
rect 46527 16544 46572 16572
rect 45235 16541 45247 16544
rect 45189 16535 45247 16541
rect 46566 16532 46572 16544
rect 46624 16532 46630 16584
rect 46676 16572 46704 16612
rect 46937 16575 46995 16581
rect 46937 16572 46949 16575
rect 46676 16544 46949 16572
rect 46937 16541 46949 16544
rect 46983 16541 46995 16575
rect 46937 16535 46995 16541
rect 48133 16575 48191 16581
rect 48133 16541 48145 16575
rect 48179 16541 48191 16575
rect 48133 16535 48191 16541
rect 40310 16504 40316 16516
rect 36096 16476 37964 16504
rect 40271 16476 40316 16504
rect 40310 16464 40316 16476
rect 40368 16464 40374 16516
rect 41230 16464 41236 16516
rect 41288 16504 41294 16516
rect 42705 16507 42763 16513
rect 42705 16504 42717 16507
rect 41288 16476 42717 16504
rect 41288 16464 41294 16476
rect 42705 16473 42717 16476
rect 42751 16504 42763 16507
rect 45002 16504 45008 16516
rect 42751 16476 45008 16504
rect 42751 16473 42763 16476
rect 42705 16467 42763 16473
rect 45002 16464 45008 16476
rect 45060 16464 45066 16516
rect 45094 16464 45100 16516
rect 45152 16504 45158 16516
rect 45152 16476 45416 16504
rect 45152 16464 45158 16476
rect 18248 16408 18552 16436
rect 18141 16399 18199 16405
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 25314 16436 25320 16448
rect 22152 16408 25320 16436
rect 22152 16396 22158 16408
rect 25314 16396 25320 16408
rect 25372 16396 25378 16448
rect 28994 16396 29000 16448
rect 29052 16436 29058 16448
rect 29917 16439 29975 16445
rect 29917 16436 29929 16439
rect 29052 16408 29929 16436
rect 29052 16396 29058 16408
rect 29917 16405 29929 16408
rect 29963 16405 29975 16439
rect 29917 16399 29975 16405
rect 30742 16396 30748 16448
rect 30800 16436 30806 16448
rect 30837 16439 30895 16445
rect 30837 16436 30849 16439
rect 30800 16408 30849 16436
rect 30800 16396 30806 16408
rect 30837 16405 30849 16408
rect 30883 16405 30895 16439
rect 33870 16436 33876 16448
rect 33831 16408 33876 16436
rect 30837 16399 30895 16405
rect 33870 16396 33876 16408
rect 33928 16396 33934 16448
rect 35437 16439 35495 16445
rect 35437 16405 35449 16439
rect 35483 16436 35495 16439
rect 35526 16436 35532 16448
rect 35483 16408 35532 16436
rect 35483 16405 35495 16408
rect 35437 16399 35495 16405
rect 35526 16396 35532 16408
rect 35584 16396 35590 16448
rect 36725 16439 36783 16445
rect 36725 16405 36737 16439
rect 36771 16436 36783 16439
rect 37274 16436 37280 16448
rect 36771 16408 37280 16436
rect 36771 16405 36783 16408
rect 36725 16399 36783 16405
rect 37274 16396 37280 16408
rect 37332 16396 37338 16448
rect 40954 16436 40960 16448
rect 40915 16408 40960 16436
rect 40954 16396 40960 16408
rect 41012 16396 41018 16448
rect 42915 16439 42973 16445
rect 42915 16405 42927 16439
rect 42961 16436 42973 16439
rect 43533 16439 43591 16445
rect 43533 16436 43545 16439
rect 42961 16408 43545 16436
rect 42961 16405 42973 16408
rect 42915 16399 42973 16405
rect 43533 16405 43545 16408
rect 43579 16405 43591 16439
rect 45278 16436 45284 16448
rect 45239 16408 45284 16436
rect 43533 16399 43591 16405
rect 45278 16396 45284 16408
rect 45336 16396 45342 16448
rect 45388 16445 45416 16476
rect 45462 16464 45468 16516
rect 45520 16504 45526 16516
rect 46845 16507 46903 16513
rect 46845 16504 46857 16507
rect 45520 16476 46857 16504
rect 45520 16464 45526 16476
rect 46845 16473 46857 16476
rect 46891 16473 46903 16507
rect 46845 16467 46903 16473
rect 47026 16464 47032 16516
rect 47084 16513 47090 16516
rect 47084 16507 47112 16513
rect 47100 16473 47112 16507
rect 48148 16504 48176 16535
rect 47084 16467 47112 16473
rect 47228 16476 48176 16504
rect 47084 16464 47090 16467
rect 47228 16445 47256 16476
rect 45373 16439 45431 16445
rect 45373 16405 45385 16439
rect 45419 16405 45431 16439
rect 45373 16399 45431 16405
rect 47213 16439 47271 16445
rect 47213 16405 47225 16439
rect 47259 16405 47271 16439
rect 47946 16436 47952 16448
rect 47907 16408 47952 16436
rect 47213 16399 47271 16405
rect 47946 16396 47952 16408
rect 48004 16396 48010 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 2406 16232 2412 16244
rect 2367 16204 2412 16232
rect 2406 16192 2412 16204
rect 2464 16192 2470 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 2832 16204 2877 16232
rect 2832 16192 2838 16204
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 6696 16204 7757 16232
rect 6696 16192 6702 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 7745 16195 7803 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 18049 16235 18107 16241
rect 18049 16232 18061 16235
rect 10928 16204 18061 16232
rect 10928 16192 10934 16204
rect 18049 16201 18061 16204
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 18380 16204 19073 16232
rect 18380 16192 18386 16204
rect 19061 16201 19073 16204
rect 19107 16201 19119 16235
rect 24946 16232 24952 16244
rect 19061 16195 19119 16201
rect 21008 16204 24952 16232
rect 2314 16124 2320 16176
rect 2372 16164 2378 16176
rect 15378 16164 15384 16176
rect 2372 16136 15384 16164
rect 2372 16124 2378 16136
rect 15378 16124 15384 16136
rect 15436 16124 15442 16176
rect 17420 16136 18460 16164
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16096 2927 16099
rect 3786 16096 3792 16108
rect 2915 16068 3792 16096
rect 2915 16065 2927 16068
rect 2869 16059 2927 16065
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 6270 16056 6276 16108
rect 6328 16096 6334 16108
rect 6621 16099 6679 16105
rect 6621 16096 6633 16099
rect 6328 16068 6633 16096
rect 6328 16056 6334 16068
rect 6621 16065 6633 16068
rect 6667 16065 6679 16099
rect 6621 16059 6679 16065
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10560 16068 10977 16096
rect 10560 16056 10566 16068
rect 10965 16065 10977 16068
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 14458 16096 14464 16108
rect 13403 16068 14464 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14636 16099 14694 16105
rect 14636 16065 14648 16099
rect 14682 16096 14694 16099
rect 14918 16096 14924 16108
rect 14682 16068 14924 16096
rect 14682 16065 14694 16068
rect 14636 16059 14694 16065
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 17420 16105 17448 16136
rect 18432 16108 18460 16136
rect 18782 16124 18788 16176
rect 18840 16164 18846 16176
rect 20717 16167 20775 16173
rect 20717 16164 20729 16167
rect 18840 16136 20729 16164
rect 18840 16124 18846 16136
rect 20717 16133 20729 16136
rect 20763 16133 20775 16167
rect 20898 16164 20904 16176
rect 20859 16136 20904 16164
rect 20717 16127 20775 16133
rect 20898 16124 20904 16136
rect 20956 16124 20962 16176
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 17494 16056 17500 16108
rect 17552 16096 17558 16108
rect 18230 16096 18236 16108
rect 17552 16068 17597 16096
rect 18191 16068 18236 16096
rect 17552 16056 17558 16068
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18414 16096 18420 16108
rect 18375 16068 18420 16096
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16096 18567 16099
rect 18690 16096 18696 16108
rect 18555 16068 18696 16096
rect 18555 16065 18567 16068
rect 18509 16059 18567 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19058 16056 19064 16108
rect 19116 16096 19122 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19116 16068 19257 16096
rect 19116 16056 19122 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16096 19487 16099
rect 21008 16096 21036 16204
rect 24946 16192 24952 16204
rect 25004 16232 25010 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 25004 16204 25329 16232
rect 25004 16192 25010 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 25317 16195 25375 16201
rect 28629 16235 28687 16241
rect 28629 16201 28641 16235
rect 28675 16201 28687 16235
rect 28629 16195 28687 16201
rect 30653 16235 30711 16241
rect 30653 16201 30665 16235
rect 30699 16232 30711 16235
rect 31110 16232 31116 16244
rect 30699 16204 31116 16232
rect 30699 16201 30711 16204
rect 30653 16195 30711 16201
rect 21634 16124 21640 16176
rect 21692 16164 21698 16176
rect 21692 16136 23980 16164
rect 21692 16124 21698 16136
rect 21836 16105 21864 16136
rect 23952 16108 23980 16136
rect 24118 16124 24124 16176
rect 24176 16164 24182 16176
rect 28644 16164 28672 16195
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 32401 16235 32459 16241
rect 32401 16232 32413 16235
rect 31726 16204 32413 16232
rect 29518 16167 29576 16173
rect 29518 16164 29530 16167
rect 24176 16136 28580 16164
rect 28644 16136 29530 16164
rect 24176 16124 24182 16136
rect 19475 16068 21036 16096
rect 21821 16099 21879 16105
rect 19475 16065 19487 16068
rect 19429 16059 19487 16065
rect 21821 16065 21833 16099
rect 21867 16065 21879 16099
rect 21821 16059 21879 16065
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22077 16099 22135 16105
rect 22077 16096 22089 16099
rect 21968 16068 22089 16096
rect 21968 16056 21974 16068
rect 22077 16065 22089 16068
rect 22123 16065 22135 16099
rect 23934 16096 23940 16108
rect 23895 16068 23940 16096
rect 22077 16059 22135 16065
rect 23934 16056 23940 16068
rect 23992 16056 23998 16108
rect 24204 16099 24262 16105
rect 24204 16065 24216 16099
rect 24250 16096 24262 16099
rect 24578 16096 24584 16108
rect 24250 16068 24584 16096
rect 24250 16065 24262 16068
rect 24204 16059 24262 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 28552 16096 28580 16136
rect 29518 16133 29530 16136
rect 29564 16133 29576 16167
rect 29518 16127 29576 16133
rect 30466 16124 30472 16176
rect 30524 16164 30530 16176
rect 31726 16164 31754 16204
rect 32401 16201 32413 16204
rect 32447 16201 32459 16235
rect 33134 16232 33140 16244
rect 33095 16204 33140 16232
rect 32401 16195 32459 16201
rect 33134 16192 33140 16204
rect 33192 16192 33198 16244
rect 41138 16232 41144 16244
rect 33428 16204 41144 16232
rect 30524 16136 31754 16164
rect 30524 16124 30530 16136
rect 32122 16124 32128 16176
rect 32180 16164 32186 16176
rect 32677 16167 32735 16173
rect 32677 16164 32689 16167
rect 32180 16136 32689 16164
rect 32180 16124 32186 16136
rect 32677 16133 32689 16136
rect 32723 16133 32735 16167
rect 32677 16127 32735 16133
rect 28626 16096 28632 16108
rect 28552 16068 28632 16096
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 28813 16099 28871 16105
rect 28813 16065 28825 16099
rect 28859 16096 28871 16099
rect 28994 16096 29000 16108
rect 28859 16068 29000 16096
rect 28859 16065 28871 16068
rect 28813 16059 28871 16065
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 29362 16056 29368 16108
rect 29420 16096 29426 16108
rect 31110 16096 31116 16108
rect 29420 16068 30328 16096
rect 31071 16068 31116 16096
rect 29420 16056 29426 16068
rect 3050 16028 3056 16040
rect 3011 16000 3056 16028
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 4856 16000 6377 16028
rect 4856 15988 4862 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 1854 15892 1860 15904
rect 1815 15864 1860 15892
rect 1854 15852 1860 15864
rect 1912 15852 1918 15904
rect 6380 15892 6408 15991
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 11882 16028 11888 16040
rect 8168 16000 11888 16028
rect 8168 15988 8174 16000
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14366 16028 14372 16040
rect 13872 16000 14372 16028
rect 13872 15988 13878 16000
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 17034 16028 17040 16040
rect 16995 16000 17040 16028
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 15746 15960 15752 15972
rect 15707 15932 15752 15960
rect 15746 15920 15752 15932
rect 15804 15920 15810 15972
rect 17236 15960 17264 15991
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 18326 16031 18384 16037
rect 17368 16000 17413 16028
rect 17368 15988 17374 16000
rect 18326 15997 18338 16031
rect 18372 16028 18384 16031
rect 18782 16028 18788 16040
rect 18372 16000 18788 16028
rect 18372 15997 18384 16000
rect 18326 15991 18384 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 19337 16031 19395 16037
rect 19337 16028 19349 16031
rect 19024 16000 19349 16028
rect 19024 15988 19030 16000
rect 19337 15997 19349 16000
rect 19383 15997 19395 16031
rect 19337 15991 19395 15997
rect 19521 16031 19579 16037
rect 19521 15997 19533 16031
rect 19567 15997 19579 16031
rect 29270 16028 29276 16040
rect 29231 16000 29276 16028
rect 19521 15991 19579 15997
rect 19150 15960 19156 15972
rect 17236 15932 19156 15960
rect 19150 15920 19156 15932
rect 19208 15920 19214 15972
rect 19536 15960 19564 15991
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 30300 16028 30328 16068
rect 31110 16056 31116 16068
rect 31168 16096 31174 16108
rect 32309 16099 32367 16105
rect 32309 16096 32321 16099
rect 31168 16068 32321 16096
rect 31168 16056 31174 16068
rect 32309 16065 32321 16068
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 33428 16105 33456 16204
rect 41138 16192 41144 16204
rect 41196 16192 41202 16244
rect 44913 16235 44971 16241
rect 44913 16201 44925 16235
rect 44959 16232 44971 16235
rect 45278 16232 45284 16244
rect 44959 16204 45284 16232
rect 44959 16201 44971 16204
rect 44913 16195 44971 16201
rect 45278 16192 45284 16204
rect 45336 16192 45342 16244
rect 46385 16235 46443 16241
rect 46385 16201 46397 16235
rect 46431 16232 46443 16235
rect 47026 16232 47032 16244
rect 46431 16204 47032 16232
rect 46431 16201 46443 16204
rect 46385 16195 46443 16201
rect 47026 16192 47032 16204
rect 47084 16192 47090 16244
rect 49697 16235 49755 16241
rect 49697 16232 49709 16235
rect 47596 16204 49709 16232
rect 34422 16173 34428 16176
rect 34416 16164 34428 16173
rect 34383 16136 34428 16164
rect 34416 16127 34428 16136
rect 34422 16124 34428 16127
rect 34480 16124 34486 16176
rect 34514 16124 34520 16176
rect 34572 16124 34578 16176
rect 40580 16167 40638 16173
rect 40580 16133 40592 16167
rect 40626 16164 40638 16167
rect 40954 16164 40960 16176
rect 40626 16136 40960 16164
rect 40626 16133 40638 16136
rect 40580 16127 40638 16133
rect 40954 16124 40960 16136
rect 41012 16124 41018 16176
rect 43806 16124 43812 16176
rect 43864 16164 43870 16176
rect 43864 16136 44772 16164
rect 43864 16124 43870 16136
rect 32493 16099 32551 16105
rect 32493 16096 32505 16099
rect 32456 16068 32505 16096
rect 32456 16056 32462 16068
rect 32493 16065 32505 16068
rect 32539 16065 32551 16099
rect 33413 16099 33471 16105
rect 33413 16096 33425 16099
rect 32493 16059 32551 16065
rect 32600 16068 33425 16096
rect 32600 16028 32628 16068
rect 33413 16065 33425 16068
rect 33459 16065 33471 16099
rect 33413 16059 33471 16065
rect 33597 16099 33655 16105
rect 33597 16065 33609 16099
rect 33643 16096 33655 16099
rect 33870 16096 33876 16108
rect 33643 16068 33876 16096
rect 33643 16065 33655 16068
rect 33597 16059 33655 16065
rect 33870 16056 33876 16068
rect 33928 16056 33934 16108
rect 34149 16099 34207 16105
rect 34149 16065 34161 16099
rect 34195 16096 34207 16099
rect 34532 16096 34560 16124
rect 34195 16068 34560 16096
rect 34195 16065 34207 16068
rect 34149 16059 34207 16065
rect 40218 16056 40224 16108
rect 40276 16096 40282 16108
rect 40313 16099 40371 16105
rect 40313 16096 40325 16099
rect 40276 16068 40325 16096
rect 40276 16056 40282 16068
rect 40313 16065 40325 16068
rect 40359 16096 40371 16099
rect 41046 16096 41052 16108
rect 40359 16068 41052 16096
rect 40359 16065 40371 16068
rect 40313 16059 40371 16065
rect 41046 16056 41052 16068
rect 41104 16056 41110 16108
rect 43714 16056 43720 16108
rect 43772 16096 43778 16108
rect 44100 16105 44128 16136
rect 44744 16105 44772 16136
rect 46216 16136 46888 16164
rect 43901 16099 43959 16105
rect 43901 16096 43913 16099
rect 43772 16068 43913 16096
rect 43772 16056 43778 16068
rect 43901 16065 43913 16068
rect 43947 16065 43959 16099
rect 43901 16059 43959 16065
rect 44085 16099 44143 16105
rect 44085 16065 44097 16099
rect 44131 16065 44143 16099
rect 44085 16059 44143 16065
rect 44545 16099 44603 16105
rect 44545 16065 44557 16099
rect 44591 16065 44603 16099
rect 44545 16059 44603 16065
rect 44729 16099 44787 16105
rect 44729 16065 44741 16099
rect 44775 16096 44787 16099
rect 45186 16096 45192 16108
rect 44775 16068 45192 16096
rect 44775 16065 44787 16068
rect 44729 16059 44787 16065
rect 33318 16028 33324 16040
rect 30300 16000 32628 16028
rect 33279 16000 33324 16028
rect 33318 15988 33324 16000
rect 33376 15988 33382 16040
rect 33505 16031 33563 16037
rect 33505 15997 33517 16031
rect 33551 16028 33563 16031
rect 33962 16028 33968 16040
rect 33551 16000 33968 16028
rect 33551 15997 33563 16000
rect 33505 15991 33563 15997
rect 19260 15932 19564 15960
rect 19260 15904 19288 15932
rect 26326 15920 26332 15972
rect 26384 15960 26390 15972
rect 27982 15960 27988 15972
rect 26384 15932 27988 15960
rect 26384 15920 26390 15932
rect 27982 15920 27988 15932
rect 28040 15920 28046 15972
rect 30208 15932 31754 15960
rect 7834 15892 7840 15904
rect 6380 15864 7840 15892
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8110 15892 8116 15904
rect 7984 15864 8116 15892
rect 7984 15852 7990 15864
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 10928 15864 13461 15892
rect 10928 15852 10934 15864
rect 13449 15861 13461 15864
rect 13495 15892 13507 15895
rect 18046 15892 18052 15904
rect 13495 15864 18052 15892
rect 13495 15861 13507 15864
rect 13449 15855 13507 15861
rect 18046 15852 18052 15864
rect 18104 15892 18110 15904
rect 18966 15892 18972 15904
rect 18104 15864 18972 15892
rect 18104 15852 18110 15864
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 19242 15852 19248 15904
rect 19300 15852 19306 15904
rect 20346 15892 20352 15904
rect 20307 15864 20352 15892
rect 20346 15852 20352 15864
rect 20404 15892 20410 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20404 15864 20913 15892
rect 20404 15852 20410 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15892 21143 15895
rect 22002 15892 22008 15904
rect 21131 15864 22008 15892
rect 21131 15861 21143 15864
rect 21085 15855 21143 15861
rect 22002 15852 22008 15864
rect 22060 15852 22066 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 23201 15895 23259 15901
rect 23201 15892 23213 15895
rect 22244 15864 23213 15892
rect 22244 15852 22250 15864
rect 23201 15861 23213 15864
rect 23247 15861 23259 15895
rect 23201 15855 23259 15861
rect 26418 15852 26424 15904
rect 26476 15892 26482 15904
rect 30208 15892 30236 15932
rect 26476 15864 30236 15892
rect 26476 15852 26482 15864
rect 30282 15852 30288 15904
rect 30340 15892 30346 15904
rect 30926 15892 30932 15904
rect 30340 15864 30932 15892
rect 30340 15852 30346 15864
rect 30926 15852 30932 15864
rect 30984 15892 30990 15904
rect 31205 15895 31263 15901
rect 31205 15892 31217 15895
rect 30984 15864 31217 15892
rect 30984 15852 30990 15864
rect 31205 15861 31217 15864
rect 31251 15861 31263 15895
rect 31726 15892 31754 15932
rect 32122 15920 32128 15972
rect 32180 15960 32186 15972
rect 33520 15960 33548 15991
rect 33962 15988 33968 16000
rect 34020 15988 34026 16040
rect 43916 16028 43944 16059
rect 44560 16028 44588 16059
rect 45186 16056 45192 16068
rect 45244 16056 45250 16108
rect 46216 16105 46244 16136
rect 46860 16105 46888 16136
rect 47596 16108 47624 16204
rect 49697 16201 49709 16204
rect 49743 16201 49755 16235
rect 49697 16195 49755 16201
rect 47946 16124 47952 16176
rect 48004 16164 48010 16176
rect 48562 16167 48620 16173
rect 48562 16164 48574 16167
rect 48004 16136 48574 16164
rect 48004 16124 48010 16136
rect 48562 16133 48574 16136
rect 48608 16133 48620 16167
rect 48562 16127 48620 16133
rect 46201 16099 46259 16105
rect 46201 16065 46213 16099
rect 46247 16065 46259 16099
rect 46201 16059 46259 16065
rect 46385 16099 46443 16105
rect 46385 16065 46397 16099
rect 46431 16065 46443 16099
rect 46385 16059 46443 16065
rect 46845 16099 46903 16105
rect 46845 16065 46857 16099
rect 46891 16096 46903 16099
rect 46934 16096 46940 16108
rect 46891 16068 46940 16096
rect 46891 16065 46903 16068
rect 46845 16059 46903 16065
rect 46400 16028 46428 16059
rect 46934 16056 46940 16068
rect 46992 16056 46998 16108
rect 47029 16099 47087 16105
rect 47029 16065 47041 16099
rect 47075 16065 47087 16099
rect 47578 16096 47584 16108
rect 47491 16068 47584 16096
rect 47029 16059 47087 16065
rect 47044 16028 47072 16059
rect 47578 16056 47584 16068
rect 47636 16056 47642 16108
rect 48317 16099 48375 16105
rect 48317 16065 48329 16099
rect 48363 16096 48375 16099
rect 48406 16096 48412 16108
rect 48363 16068 48412 16096
rect 48363 16065 48375 16068
rect 48317 16059 48375 16065
rect 48406 16056 48412 16068
rect 48464 16056 48470 16108
rect 47673 16031 47731 16037
rect 47673 16028 47685 16031
rect 43916 16000 45324 16028
rect 46400 16000 47685 16028
rect 32180 15932 32225 15960
rect 32692 15932 33548 15960
rect 45296 15960 45324 16000
rect 47673 15997 47685 16000
rect 47719 15997 47731 16031
rect 47673 15991 47731 15997
rect 46566 15960 46572 15972
rect 45296 15932 46572 15960
rect 32180 15920 32186 15932
rect 32692 15892 32720 15932
rect 46566 15920 46572 15932
rect 46624 15960 46630 15972
rect 46845 15963 46903 15969
rect 46845 15960 46857 15963
rect 46624 15932 46857 15960
rect 46624 15920 46630 15932
rect 46845 15929 46857 15932
rect 46891 15929 46903 15963
rect 46845 15923 46903 15929
rect 31726 15864 32720 15892
rect 31205 15855 31263 15861
rect 33502 15852 33508 15904
rect 33560 15892 33566 15904
rect 35529 15895 35587 15901
rect 35529 15892 35541 15895
rect 33560 15864 35541 15892
rect 33560 15852 33566 15864
rect 35529 15861 35541 15864
rect 35575 15861 35587 15895
rect 41690 15892 41696 15904
rect 41651 15864 41696 15892
rect 35529 15855 35587 15861
rect 41690 15852 41696 15864
rect 41748 15852 41754 15904
rect 41966 15852 41972 15904
rect 42024 15892 42030 15904
rect 43993 15895 44051 15901
rect 43993 15892 44005 15895
rect 42024 15864 44005 15892
rect 42024 15852 42030 15864
rect 43993 15861 44005 15864
rect 44039 15892 44051 15895
rect 45094 15892 45100 15904
rect 44039 15864 45100 15892
rect 44039 15861 44051 15864
rect 43993 15855 44051 15861
rect 45094 15852 45100 15864
rect 45152 15852 45158 15904
rect 45186 15852 45192 15904
rect 45244 15892 45250 15904
rect 47118 15892 47124 15904
rect 45244 15864 47124 15892
rect 45244 15852 45250 15864
rect 47118 15852 47124 15864
rect 47176 15852 47182 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2130 15648 2136 15700
rect 2188 15688 2194 15700
rect 6270 15688 6276 15700
rect 2188 15660 5957 15688
rect 6231 15660 6276 15688
rect 2188 15648 2194 15660
rect 2225 15623 2283 15629
rect 2225 15589 2237 15623
rect 2271 15620 2283 15623
rect 2866 15620 2872 15632
rect 2271 15592 2872 15620
rect 2271 15589 2283 15592
rect 2225 15583 2283 15589
rect 2866 15580 2872 15592
rect 2924 15580 2930 15632
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 3050 15552 3056 15564
rect 2823 15524 3056 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 3510 15484 3516 15496
rect 2639 15456 3516 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 1412 15416 1440 15447
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 3970 15484 3976 15496
rect 3931 15456 3976 15484
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 5626 15416 5632 15428
rect 1412 15388 5632 15416
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 5929 15416 5957 15660
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 10502 15688 10508 15700
rect 10463 15660 10508 15688
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 14918 15688 14924 15700
rect 14879 15660 14924 15688
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 16114 15688 16120 15700
rect 16075 15660 16120 15688
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 17954 15688 17960 15700
rect 16224 15660 17960 15688
rect 16224 15620 16252 15660
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 18230 15688 18236 15700
rect 18187 15660 18236 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 19058 15688 19064 15700
rect 18380 15660 19064 15688
rect 18380 15648 18386 15660
rect 19058 15648 19064 15660
rect 19116 15648 19122 15700
rect 19150 15648 19156 15700
rect 19208 15688 19214 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 19208 15660 19257 15688
rect 19208 15648 19214 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 24118 15688 24124 15700
rect 19245 15651 19303 15657
rect 20180 15660 24124 15688
rect 6472 15592 16252 15620
rect 16301 15623 16359 15629
rect 6472 15493 6500 15592
rect 16301 15589 16313 15623
rect 16347 15589 16359 15623
rect 16301 15583 16359 15589
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 11057 15555 11115 15561
rect 11057 15552 11069 15555
rect 10652 15524 11069 15552
rect 10652 15512 10658 15524
rect 11057 15521 11069 15524
rect 11103 15521 11115 15555
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 11057 15515 11115 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15381 15555 15439 15561
rect 15381 15521 15393 15555
rect 15427 15552 15439 15555
rect 16316 15552 16344 15583
rect 18782 15580 18788 15632
rect 18840 15620 18846 15632
rect 20180 15620 20208 15660
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24578 15688 24584 15700
rect 24539 15660 24584 15688
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 26418 15688 26424 15700
rect 24688 15660 26424 15688
rect 18840 15592 20208 15620
rect 18840 15580 18846 15592
rect 20254 15580 20260 15632
rect 20312 15620 20318 15632
rect 24688 15620 24716 15660
rect 26418 15648 26424 15660
rect 26476 15648 26482 15700
rect 26513 15691 26571 15697
rect 26513 15657 26525 15691
rect 26559 15688 26571 15691
rect 26602 15688 26608 15700
rect 26559 15660 26608 15688
rect 26559 15657 26571 15660
rect 26513 15651 26571 15657
rect 26602 15648 26608 15660
rect 26660 15688 26666 15700
rect 26660 15660 28994 15688
rect 26660 15648 26666 15660
rect 26697 15623 26755 15629
rect 26697 15620 26709 15623
rect 20312 15592 24716 15620
rect 24780 15592 26709 15620
rect 20312 15580 20318 15592
rect 15427 15524 16344 15552
rect 15427 15521 15439 15524
rect 15381 15515 15439 15521
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 18417 15555 18475 15561
rect 18417 15552 18429 15555
rect 18104 15524 18429 15552
rect 18104 15512 18110 15524
rect 18417 15521 18429 15524
rect 18463 15521 18475 15555
rect 18598 15552 18604 15564
rect 18559 15524 18604 15552
rect 18417 15515 18475 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 19058 15512 19064 15564
rect 19116 15552 19122 15564
rect 19429 15555 19487 15561
rect 19429 15552 19441 15555
rect 19116 15524 19441 15552
rect 19116 15512 19122 15524
rect 19429 15521 19441 15524
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15552 19671 15555
rect 19659 15524 22232 15552
rect 19659 15521 19671 15524
rect 19613 15515 19671 15521
rect 22204 15496 22232 15524
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6638 15484 6644 15496
rect 6599 15456 6644 15484
rect 6457 15447 6515 15453
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 10870 15484 10876 15496
rect 6788 15456 6833 15484
rect 10831 15456 10876 15484
rect 6788 15444 6794 15456
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 18322 15484 18328 15496
rect 18283 15456 18328 15484
rect 15197 15447 15255 15453
rect 15212 15416 15240 15447
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 18564 15456 18609 15484
rect 18564 15444 18570 15456
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19024 15456 19533 15484
rect 19024 15444 19030 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 22002 15484 22008 15496
rect 21963 15456 22008 15484
rect 19705 15447 19763 15453
rect 15378 15416 15384 15428
rect 5929 15388 12434 15416
rect 15212 15388 15384 15416
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 2685 15351 2743 15357
rect 2685 15317 2697 15351
rect 2731 15348 2743 15351
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 2731 15320 3801 15348
rect 2731 15317 2743 15320
rect 2685 15311 2743 15317
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3789 15311 3847 15317
rect 10965 15351 11023 15357
rect 10965 15317 10977 15351
rect 11011 15348 11023 15351
rect 11054 15348 11060 15360
rect 11011 15320 11060 15348
rect 11011 15317 11023 15320
rect 10965 15311 11023 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12406 15348 12434 15388
rect 15378 15376 15384 15388
rect 15436 15376 15442 15428
rect 15746 15376 15752 15428
rect 15804 15416 15810 15428
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 15804 15388 15945 15416
rect 15804 15376 15810 15388
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 15933 15379 15991 15385
rect 16040 15388 18552 15416
rect 16040 15348 16068 15388
rect 12406 15320 16068 15348
rect 16143 15351 16201 15357
rect 16143 15317 16155 15351
rect 16189 15348 16201 15351
rect 16298 15348 16304 15360
rect 16189 15320 16304 15348
rect 16189 15317 16201 15320
rect 16143 15311 16201 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 18524 15348 18552 15388
rect 18598 15376 18604 15428
rect 18656 15416 18662 15428
rect 19242 15416 19248 15428
rect 18656 15388 19248 15416
rect 18656 15376 18662 15388
rect 19242 15376 19248 15388
rect 19300 15416 19306 15428
rect 19720 15416 19748 15447
rect 22002 15444 22008 15456
rect 22060 15484 22066 15496
rect 22186 15484 22192 15496
rect 22060 15444 22094 15484
rect 22147 15456 22192 15484
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15484 22339 15487
rect 22646 15484 22652 15496
rect 22327 15456 22652 15484
rect 22327 15453 22339 15456
rect 22281 15447 22339 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 24780 15493 24808 15592
rect 26697 15589 26709 15592
rect 26743 15589 26755 15623
rect 26697 15583 26755 15589
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25961 15555 26019 15561
rect 25961 15552 25973 15555
rect 24912 15524 25973 15552
rect 24912 15512 24918 15524
rect 25961 15521 25973 15524
rect 26007 15552 26019 15555
rect 26602 15552 26608 15564
rect 26007 15524 26608 15552
rect 26007 15521 26019 15524
rect 25961 15515 26019 15521
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24946 15484 24952 15496
rect 24907 15456 24952 15484
rect 24765 15447 24823 15453
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 25041 15487 25099 15493
rect 25041 15453 25053 15487
rect 25087 15484 25099 15487
rect 25406 15484 25412 15496
rect 25087 15456 25412 15484
rect 25087 15453 25099 15456
rect 25041 15447 25099 15453
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 26712 15484 26740 15583
rect 28966 15552 28994 15660
rect 29546 15648 29552 15700
rect 29604 15688 29610 15700
rect 30285 15691 30343 15697
rect 30285 15688 30297 15691
rect 29604 15660 30297 15688
rect 29604 15648 29610 15660
rect 30285 15657 30297 15660
rect 30331 15657 30343 15691
rect 33597 15691 33655 15697
rect 33597 15688 33609 15691
rect 30285 15651 30343 15657
rect 31726 15660 33609 15688
rect 30193 15623 30251 15629
rect 30193 15589 30205 15623
rect 30239 15620 30251 15623
rect 30742 15620 30748 15632
rect 30239 15592 30748 15620
rect 30239 15589 30251 15592
rect 30193 15583 30251 15589
rect 30742 15580 30748 15592
rect 30800 15620 30806 15632
rect 31726 15620 31754 15660
rect 33597 15657 33609 15660
rect 33643 15657 33655 15691
rect 33597 15651 33655 15657
rect 33689 15691 33747 15697
rect 33689 15657 33701 15691
rect 33735 15688 33747 15691
rect 33778 15688 33784 15700
rect 33735 15660 33784 15688
rect 33735 15657 33747 15660
rect 33689 15651 33747 15657
rect 33778 15648 33784 15660
rect 33836 15648 33842 15700
rect 33962 15648 33968 15700
rect 34020 15688 34026 15700
rect 35069 15691 35127 15697
rect 35069 15688 35081 15691
rect 34020 15660 35081 15688
rect 34020 15648 34026 15660
rect 35069 15657 35081 15660
rect 35115 15657 35127 15691
rect 40586 15688 40592 15700
rect 35069 15651 35127 15657
rect 35176 15660 40264 15688
rect 40547 15660 40592 15688
rect 30800 15592 31754 15620
rect 30800 15580 30806 15592
rect 32766 15580 32772 15632
rect 32824 15620 32830 15632
rect 35176 15620 35204 15660
rect 36262 15620 36268 15632
rect 32824 15592 35204 15620
rect 35268 15592 36268 15620
rect 32824 15580 32830 15592
rect 33781 15555 33839 15561
rect 28966 15524 33640 15552
rect 27341 15487 27399 15493
rect 27341 15484 27353 15487
rect 25884 15456 26648 15484
rect 26712 15456 27353 15484
rect 19300 15388 19748 15416
rect 21821 15419 21879 15425
rect 19300 15376 19306 15388
rect 21821 15385 21833 15419
rect 21867 15416 21879 15419
rect 21910 15416 21916 15428
rect 21867 15388 21916 15416
rect 21867 15385 21879 15388
rect 21821 15379 21879 15385
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 20346 15348 20352 15360
rect 18524 15320 20352 15348
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 22066 15348 22094 15444
rect 25884 15348 25912 15456
rect 26326 15416 26332 15428
rect 26287 15388 26332 15416
rect 26326 15376 26332 15388
rect 26384 15376 26390 15428
rect 26510 15376 26516 15428
rect 26568 15425 26574 15428
rect 26568 15419 26587 15425
rect 26575 15385 26587 15419
rect 26568 15379 26587 15385
rect 26568 15376 26574 15379
rect 22066 15320 25912 15348
rect 26620 15348 26648 15456
rect 27341 15453 27353 15456
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 30101 15487 30159 15493
rect 30101 15453 30113 15487
rect 30147 15484 30159 15487
rect 30190 15484 30196 15496
rect 30147 15456 30196 15484
rect 30147 15453 30159 15456
rect 30101 15447 30159 15453
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30282 15444 30288 15496
rect 30340 15484 30346 15496
rect 30558 15484 30564 15496
rect 30340 15456 30564 15484
rect 30340 15444 30346 15456
rect 30558 15444 30564 15456
rect 30616 15444 30622 15496
rect 32122 15444 32128 15496
rect 32180 15484 32186 15496
rect 33502 15484 33508 15496
rect 32180 15456 33508 15484
rect 32180 15444 32186 15456
rect 33502 15444 33508 15456
rect 33560 15444 33566 15496
rect 33612 15484 33640 15524
rect 33781 15521 33793 15555
rect 33827 15552 33839 15555
rect 34054 15552 34060 15564
rect 33827 15524 34060 15552
rect 33827 15521 33839 15524
rect 33781 15515 33839 15521
rect 34054 15512 34060 15524
rect 34112 15512 34118 15564
rect 35268 15552 35296 15592
rect 36262 15580 36268 15592
rect 36320 15580 36326 15632
rect 37366 15580 37372 15632
rect 37424 15620 37430 15632
rect 37645 15623 37703 15629
rect 37645 15620 37657 15623
rect 37424 15592 37657 15620
rect 37424 15580 37430 15592
rect 37645 15589 37657 15592
rect 37691 15589 37703 15623
rect 37645 15583 37703 15589
rect 34164 15524 35296 15552
rect 35713 15555 35771 15561
rect 34164 15484 34192 15524
rect 35713 15521 35725 15555
rect 35759 15552 35771 15555
rect 38654 15552 38660 15564
rect 35759 15524 38660 15552
rect 35759 15521 35771 15524
rect 35713 15515 35771 15521
rect 33612 15456 34192 15484
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34848 15456 34897 15484
rect 34848 15444 34854 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 27154 15416 27160 15428
rect 27115 15388 27160 15416
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 29917 15419 29975 15425
rect 27448 15388 29868 15416
rect 27448 15348 27476 15388
rect 26620 15320 27476 15348
rect 27525 15351 27583 15357
rect 27525 15317 27537 15351
rect 27571 15348 27583 15351
rect 28258 15348 28264 15360
rect 27571 15320 28264 15348
rect 27571 15317 27583 15320
rect 27525 15311 27583 15317
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 29840 15348 29868 15388
rect 29917 15385 29929 15419
rect 29963 15416 29975 15419
rect 30374 15416 30380 15428
rect 29963 15388 30380 15416
rect 29963 15385 29975 15388
rect 29917 15379 29975 15385
rect 30374 15376 30380 15388
rect 30432 15376 30438 15428
rect 31294 15376 31300 15428
rect 31352 15416 31358 15428
rect 31478 15416 31484 15428
rect 31352 15388 31484 15416
rect 31352 15376 31358 15388
rect 31478 15376 31484 15388
rect 31536 15376 31542 15428
rect 31018 15348 31024 15360
rect 29840 15320 31024 15348
rect 31018 15308 31024 15320
rect 31076 15308 31082 15360
rect 31202 15308 31208 15360
rect 31260 15348 31266 15360
rect 35728 15348 35756 15515
rect 38654 15512 38660 15524
rect 38712 15512 38718 15564
rect 40236 15561 40264 15660
rect 40586 15648 40592 15660
rect 40644 15648 40650 15700
rect 54754 15688 54760 15700
rect 54715 15660 54760 15688
rect 54754 15648 54760 15660
rect 54812 15648 54818 15700
rect 41690 15580 41696 15632
rect 41748 15620 41754 15632
rect 41748 15592 42196 15620
rect 41748 15580 41754 15592
rect 40221 15555 40279 15561
rect 40221 15521 40233 15555
rect 40267 15521 40279 15555
rect 41785 15555 41843 15561
rect 41785 15552 41797 15555
rect 40221 15515 40279 15521
rect 40420 15524 41797 15552
rect 35986 15484 35992 15496
rect 35947 15456 35992 15484
rect 35986 15444 35992 15456
rect 36044 15444 36050 15496
rect 37918 15484 37924 15496
rect 37879 15456 37924 15484
rect 37918 15444 37924 15456
rect 37976 15444 37982 15496
rect 40420 15493 40448 15524
rect 41785 15521 41797 15524
rect 41831 15521 41843 15555
rect 41966 15552 41972 15564
rect 41927 15524 41972 15552
rect 41785 15515 41843 15521
rect 41966 15512 41972 15524
rect 42024 15512 42030 15564
rect 42168 15561 42196 15592
rect 42153 15555 42211 15561
rect 42153 15521 42165 15555
rect 42199 15552 42211 15555
rect 43254 15552 43260 15564
rect 42199 15524 43260 15552
rect 42199 15521 42211 15524
rect 42153 15515 42211 15521
rect 43254 15512 43260 15524
rect 43312 15552 43318 15564
rect 47578 15552 47584 15564
rect 43312 15524 43576 15552
rect 43312 15512 43318 15524
rect 40405 15487 40463 15493
rect 40405 15453 40417 15487
rect 40451 15453 40463 15487
rect 40405 15447 40463 15453
rect 40862 15444 40868 15496
rect 40920 15484 40926 15496
rect 42061 15487 42119 15493
rect 42061 15484 42073 15487
rect 40920 15456 42073 15484
rect 40920 15444 40926 15456
rect 42061 15453 42073 15456
rect 42107 15453 42119 15487
rect 42061 15447 42119 15453
rect 42245 15487 42303 15493
rect 42245 15453 42257 15487
rect 42291 15484 42303 15487
rect 43438 15484 43444 15496
rect 42291 15456 43444 15484
rect 42291 15453 42303 15456
rect 42245 15447 42303 15453
rect 43438 15444 43444 15456
rect 43496 15444 43502 15496
rect 43548 15493 43576 15524
rect 47044 15524 47584 15552
rect 43533 15487 43591 15493
rect 43533 15453 43545 15487
rect 43579 15453 43591 15487
rect 43533 15447 43591 15453
rect 43717 15487 43775 15493
rect 43717 15453 43729 15487
rect 43763 15484 43775 15487
rect 43990 15484 43996 15496
rect 43763 15456 43996 15484
rect 43763 15453 43775 15456
rect 43717 15447 43775 15453
rect 43990 15444 43996 15456
rect 44048 15444 44054 15496
rect 47044 15493 47072 15524
rect 47578 15512 47584 15524
rect 47636 15512 47642 15564
rect 47029 15487 47087 15493
rect 47029 15453 47041 15487
rect 47075 15453 47087 15487
rect 47029 15447 47087 15453
rect 47118 15444 47124 15496
rect 47176 15484 47182 15496
rect 47176 15456 47221 15484
rect 47176 15444 47182 15456
rect 53098 15444 53104 15496
rect 53156 15484 53162 15496
rect 53377 15487 53435 15493
rect 53377 15484 53389 15487
rect 53156 15456 53389 15484
rect 53156 15444 53162 15456
rect 53377 15453 53389 15456
rect 53423 15453 53435 15487
rect 53377 15447 53435 15453
rect 37642 15416 37648 15428
rect 37603 15388 37648 15416
rect 37642 15376 37648 15388
rect 37700 15376 37706 15428
rect 46845 15419 46903 15425
rect 46845 15385 46857 15419
rect 46891 15416 46903 15419
rect 47946 15416 47952 15428
rect 46891 15388 47952 15416
rect 46891 15385 46903 15388
rect 46845 15379 46903 15385
rect 47946 15376 47952 15388
rect 48004 15376 48010 15428
rect 53006 15376 53012 15428
rect 53064 15416 53070 15428
rect 53622 15419 53680 15425
rect 53622 15416 53634 15419
rect 53064 15388 53634 15416
rect 53064 15376 53070 15388
rect 53622 15385 53634 15388
rect 53668 15385 53680 15419
rect 53622 15379 53680 15385
rect 37826 15348 37832 15360
rect 31260 15320 35756 15348
rect 37739 15320 37832 15348
rect 31260 15308 31266 15320
rect 37826 15308 37832 15320
rect 37884 15348 37890 15360
rect 41230 15348 41236 15360
rect 37884 15320 41236 15348
rect 37884 15308 37890 15320
rect 41230 15308 41236 15320
rect 41288 15308 41294 15360
rect 43717 15351 43775 15357
rect 43717 15317 43729 15351
rect 43763 15348 43775 15351
rect 44358 15348 44364 15360
rect 43763 15320 44364 15348
rect 43763 15317 43775 15320
rect 43717 15311 43775 15317
rect 44358 15308 44364 15320
rect 44416 15308 44422 15360
rect 46934 15348 46940 15360
rect 46895 15320 46940 15348
rect 46934 15308 46940 15320
rect 46992 15308 46998 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1946 15144 1952 15156
rect 1859 15116 1952 15144
rect 1946 15104 1952 15116
rect 2004 15144 2010 15156
rect 4246 15144 4252 15156
rect 2004 15116 4252 15144
rect 2004 15104 2010 15116
rect 4246 15104 4252 15116
rect 4304 15144 4310 15156
rect 4798 15144 4804 15156
rect 4304 15116 4804 15144
rect 4304 15104 4310 15116
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5626 15144 5632 15156
rect 5587 15116 5632 15144
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 8202 15104 8208 15156
rect 8260 15144 8266 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 8260 15116 8677 15144
rect 8260 15104 8266 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8665 15107 8723 15113
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 9490 15144 9496 15156
rect 8803 15116 9496 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 12066 15144 12072 15156
rect 12027 15116 12072 15144
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12216 15116 17264 15144
rect 12216 15104 12222 15116
rect 1964 15017 1992 15104
rect 2590 15036 2596 15088
rect 2648 15076 2654 15088
rect 13449 15079 13507 15085
rect 2648 15048 13308 15076
rect 2648 15036 2654 15048
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 14977 2007 15011
rect 1949 14971 2007 14977
rect 2216 15011 2274 15017
rect 2216 14977 2228 15011
rect 2262 15008 2274 15011
rect 2682 15008 2688 15020
rect 2262 14980 2688 15008
rect 2262 14977 2274 14980
rect 2216 14971 2274 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 4246 15008 4252 15020
rect 3844 14980 4252 15008
rect 3844 14968 3850 14980
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4516 15011 4574 15017
rect 4516 14977 4528 15011
rect 4562 15008 4574 15011
rect 5074 15008 5080 15020
rect 4562 14980 5080 15008
rect 4562 14977 4574 14980
rect 4516 14971 4574 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7558 15008 7564 15020
rect 7423 14980 7564 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 11977 15011 12035 15017
rect 8904 14980 8949 15008
rect 8904 14968 8910 14980
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12618 15008 12624 15020
rect 12023 14980 12434 15008
rect 12579 14980 12624 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12406 14952 12434 14980
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 7064 14912 7205 14940
rect 7064 14900 7070 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8297 14943 8355 14949
rect 8297 14909 8309 14943
rect 8343 14940 8355 14943
rect 12158 14940 12164 14952
rect 8343 14912 12164 14940
rect 8343 14909 8355 14912
rect 8297 14903 8355 14909
rect 8128 14872 8156 14903
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12406 14912 12440 14952
rect 12434 14900 12440 14912
rect 12492 14940 12498 14952
rect 12820 14940 12848 14971
rect 12492 14912 12848 14940
rect 13280 14940 13308 15048
rect 13449 15045 13461 15079
rect 13495 15076 13507 15079
rect 13538 15076 13544 15088
rect 13495 15048 13544 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 13633 15079 13691 15085
rect 13633 15045 13645 15079
rect 13679 15045 13691 15079
rect 17236 15076 17264 15116
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18049 15147 18107 15153
rect 18049 15144 18061 15147
rect 18012 15116 18061 15144
rect 18012 15104 18018 15116
rect 18049 15113 18061 15116
rect 18095 15113 18107 15147
rect 18049 15107 18107 15113
rect 21818 15104 21824 15156
rect 21876 15104 21882 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22833 15147 22891 15153
rect 22833 15144 22845 15147
rect 22152 15116 22845 15144
rect 22152 15104 22158 15116
rect 22833 15113 22845 15116
rect 22879 15113 22891 15147
rect 22833 15107 22891 15113
rect 26973 15147 27031 15153
rect 26973 15113 26985 15147
rect 27019 15144 27031 15147
rect 27154 15144 27160 15156
rect 27019 15116 27160 15144
rect 27019 15113 27031 15116
rect 26973 15107 27031 15113
rect 27154 15104 27160 15116
rect 27212 15104 27218 15156
rect 30374 15104 30380 15156
rect 30432 15144 30438 15156
rect 31481 15147 31539 15153
rect 31481 15144 31493 15147
rect 30432 15116 31493 15144
rect 30432 15104 30438 15116
rect 31481 15113 31493 15116
rect 31527 15113 31539 15147
rect 31481 15107 31539 15113
rect 36722 15104 36728 15156
rect 36780 15144 36786 15156
rect 37642 15144 37648 15156
rect 36780 15116 37648 15144
rect 36780 15104 36786 15116
rect 37642 15104 37648 15116
rect 37700 15144 37706 15156
rect 38749 15147 38807 15153
rect 38749 15144 38761 15147
rect 37700 15116 38761 15144
rect 37700 15104 37706 15116
rect 38749 15113 38761 15116
rect 38795 15113 38807 15147
rect 38749 15107 38807 15113
rect 40957 15147 41015 15153
rect 40957 15113 40969 15147
rect 41003 15144 41015 15147
rect 41230 15144 41236 15156
rect 41003 15116 41236 15144
rect 41003 15113 41015 15116
rect 40957 15107 41015 15113
rect 41230 15104 41236 15116
rect 41288 15104 41294 15156
rect 43625 15147 43683 15153
rect 43625 15113 43637 15147
rect 43671 15144 43683 15147
rect 44269 15147 44327 15153
rect 44269 15144 44281 15147
rect 43671 15116 44281 15144
rect 43671 15113 43683 15116
rect 43625 15107 43683 15113
rect 44269 15113 44281 15116
rect 44315 15113 44327 15147
rect 44269 15107 44327 15113
rect 47026 15104 47032 15156
rect 47084 15144 47090 15156
rect 47673 15147 47731 15153
rect 47673 15144 47685 15147
rect 47084 15116 47685 15144
rect 47084 15104 47090 15116
rect 47673 15113 47685 15116
rect 47719 15113 47731 15147
rect 53006 15144 53012 15156
rect 52967 15116 53012 15144
rect 47673 15107 47731 15113
rect 53006 15104 53012 15116
rect 53064 15104 53070 15156
rect 21634 15076 21640 15088
rect 17236 15048 21640 15076
rect 13633 15039 13691 15045
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13648 15008 13676 15039
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 13412 14980 13676 15008
rect 14660 14980 15301 15008
rect 13412 14968 13418 14980
rect 14660 14949 14688 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 16574 15008 16580 15020
rect 15519 14980 16580 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 13280 14912 14657 14940
rect 12492 14900 12498 14912
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 15194 14940 15200 14952
rect 15155 14912 15200 14940
rect 14645 14903 14703 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 8570 14872 8576 14884
rect 8128 14844 8576 14872
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 15304 14872 15332 14971
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 15008 18567 15011
rect 18690 15008 18696 15020
rect 18555 14980 18696 15008
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20956 14980 21005 15008
rect 20956 14968 20962 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15436 14912 15481 14940
rect 15436 14900 15442 14912
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 18196 14912 18245 14940
rect 18196 14900 18202 14912
rect 18233 14909 18245 14912
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18380 14912 18425 14940
rect 18380 14900 18386 14912
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 21634 14940 21640 14952
rect 18840 14912 21640 14940
rect 18840 14900 18846 14912
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 21836 14940 21864 15104
rect 30926 15076 30932 15088
rect 27337 15048 30932 15076
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21933 14980 22017 15008
rect 21933 14940 21961 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22152 14980 22197 15008
rect 22152 14968 22158 14980
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22520 14980 22569 15008
rect 22520 14968 22526 14980
rect 22557 14977 22569 14980
rect 22603 15008 22615 15011
rect 23290 15008 23296 15020
rect 22603 14980 23296 15008
rect 22603 14977 22615 14980
rect 22557 14971 22615 14977
rect 23290 14968 23296 14980
rect 23348 14968 23354 15020
rect 27062 14968 27068 15020
rect 27120 15008 27126 15020
rect 27337 15017 27365 15048
rect 30926 15036 30932 15048
rect 30984 15036 30990 15088
rect 32398 15076 32404 15088
rect 31496 15048 32404 15076
rect 27203 15011 27261 15017
rect 27203 15008 27215 15011
rect 27120 14980 27215 15008
rect 27120 14968 27126 14980
rect 27203 14977 27215 14980
rect 27249 14977 27261 15011
rect 27203 14971 27261 14977
rect 27322 15011 27380 15017
rect 27322 14977 27334 15011
rect 27368 14977 27380 15011
rect 27322 14971 27380 14977
rect 21836 14912 21961 14940
rect 26602 14900 26608 14952
rect 26660 14940 26666 14952
rect 27337 14940 27365 14971
rect 27430 14968 27436 15020
rect 27488 15017 27494 15020
rect 27488 15008 27496 15017
rect 27488 14980 27533 15008
rect 27488 14971 27496 14980
rect 27488 14968 27494 14971
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 28258 15008 28264 15020
rect 27672 14980 27717 15008
rect 28219 14980 28264 15008
rect 27672 14968 27678 14980
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 30745 15011 30803 15017
rect 30745 15008 30757 15011
rect 30524 14980 30757 15008
rect 30524 14968 30530 14980
rect 30745 14977 30757 14980
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 15008 31447 15011
rect 31496 15008 31524 15048
rect 32398 15036 32404 15048
rect 32456 15036 32462 15088
rect 34514 15036 34520 15088
rect 34572 15076 34578 15088
rect 37274 15076 37280 15088
rect 34572 15048 37280 15076
rect 34572 15036 34578 15048
rect 37274 15036 37280 15048
rect 37332 15076 37338 15088
rect 40862 15076 40868 15088
rect 37332 15048 37412 15076
rect 40823 15048 40868 15076
rect 37332 15036 37338 15048
rect 31435 14980 31524 15008
rect 31573 15011 31631 15017
rect 31435 14977 31447 14980
rect 31389 14971 31447 14977
rect 31573 14977 31585 15011
rect 31619 14977 31631 15011
rect 31573 14971 31631 14977
rect 34425 15011 34483 15017
rect 34425 14977 34437 15011
rect 34471 15008 34483 15011
rect 35986 15008 35992 15020
rect 34471 14980 35992 15008
rect 34471 14977 34483 14980
rect 34425 14971 34483 14977
rect 26660 14912 27365 14940
rect 26660 14900 26666 14912
rect 30926 14900 30932 14952
rect 30984 14940 30990 14952
rect 31588 14940 31616 14971
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 37384 15017 37412 15048
rect 40862 15036 40868 15048
rect 40920 15036 40926 15088
rect 43714 15036 43720 15088
rect 43772 15076 43778 15088
rect 44085 15079 44143 15085
rect 44085 15076 44097 15079
rect 43772 15048 44097 15076
rect 43772 15036 43778 15048
rect 44085 15045 44097 15048
rect 44131 15076 44143 15079
rect 46934 15076 46940 15088
rect 44131 15048 46940 15076
rect 44131 15045 44143 15048
rect 44085 15039 44143 15045
rect 46934 15036 46940 15048
rect 46992 15036 46998 15088
rect 37369 15011 37427 15017
rect 37369 14977 37381 15011
rect 37415 14977 37427 15011
rect 37369 14971 37427 14977
rect 37458 14968 37464 15020
rect 37516 15008 37522 15020
rect 37625 15011 37683 15017
rect 37625 15008 37637 15011
rect 37516 14980 37637 15008
rect 37516 14968 37522 14980
rect 37625 14977 37637 14980
rect 37671 14977 37683 15011
rect 37625 14971 37683 14977
rect 38746 14968 38752 15020
rect 38804 15008 38810 15020
rect 43257 15011 43315 15017
rect 43257 15008 43269 15011
rect 38804 14980 43269 15008
rect 38804 14968 38810 14980
rect 43257 14977 43269 14980
rect 43303 14977 43315 15011
rect 43257 14971 43315 14977
rect 43441 15011 43499 15017
rect 43441 14977 43453 15011
rect 43487 15008 43499 15011
rect 43990 15008 43996 15020
rect 43487 14980 43996 15008
rect 43487 14977 43499 14980
rect 43441 14971 43499 14977
rect 43990 14968 43996 14980
rect 44048 14968 44054 15020
rect 44358 15008 44364 15020
rect 44319 14980 44364 15008
rect 44358 14968 44364 14980
rect 44416 14968 44422 15020
rect 46658 14968 46664 15020
rect 46716 15008 46722 15020
rect 47581 15011 47639 15017
rect 47581 15008 47593 15011
rect 46716 14980 47593 15008
rect 46716 14968 46722 14980
rect 47581 14977 47593 14980
rect 47627 14977 47639 15011
rect 47581 14971 47639 14977
rect 47765 15011 47823 15017
rect 47765 14977 47777 15011
rect 47811 15008 47823 15011
rect 47946 15008 47952 15020
rect 47811 14980 47952 15008
rect 47811 14977 47823 14980
rect 47765 14971 47823 14977
rect 47946 14968 47952 14980
rect 48004 14968 48010 15020
rect 53190 15008 53196 15020
rect 53151 14980 53196 15008
rect 53190 14968 53196 14980
rect 53248 14968 53254 15020
rect 30984 14912 31616 14940
rect 30984 14900 30990 14912
rect 31754 14900 31760 14952
rect 31812 14940 31818 14952
rect 36998 14940 37004 14952
rect 31812 14912 37004 14940
rect 31812 14900 31818 14912
rect 36998 14900 37004 14912
rect 37056 14900 37062 14952
rect 10192 14844 13676 14872
rect 15304 14844 22094 14872
rect 10192 14832 10198 14844
rect 3329 14807 3387 14813
rect 3329 14773 3341 14807
rect 3375 14804 3387 14807
rect 3510 14804 3516 14816
rect 3375 14776 3516 14804
rect 3375 14773 3387 14776
rect 3329 14767 3387 14773
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 7558 14804 7564 14816
rect 7519 14776 7564 14804
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 11146 14804 11152 14816
rect 10008 14776 11152 14804
rect 10008 14764 10014 14776
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 12621 14807 12679 14813
rect 12621 14773 12633 14807
rect 12667 14804 12679 14807
rect 13262 14804 13268 14816
rect 12667 14776 13268 14804
rect 12667 14773 12679 14776
rect 12621 14767 12679 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13648 14813 13676 14844
rect 13633 14807 13691 14813
rect 13633 14773 13645 14807
rect 13679 14773 13691 14807
rect 13814 14804 13820 14816
rect 13775 14776 13820 14804
rect 13633 14767 13691 14773
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 15010 14804 15016 14816
rect 14971 14776 15016 14804
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 18782 14804 18788 14816
rect 15252 14776 18788 14804
rect 15252 14764 15258 14776
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 21177 14807 21235 14813
rect 21177 14773 21189 14807
rect 21223 14804 21235 14807
rect 21634 14804 21640 14816
rect 21223 14776 21640 14804
rect 21223 14773 21235 14776
rect 21177 14767 21235 14773
rect 21634 14764 21640 14776
rect 21692 14764 21698 14816
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22066 14804 22094 14844
rect 22278 14832 22284 14884
rect 22336 14872 22342 14884
rect 32306 14872 32312 14884
rect 22336 14844 32312 14872
rect 22336 14832 22342 14844
rect 32306 14832 32312 14844
rect 32364 14832 32370 14884
rect 27890 14804 27896 14816
rect 22066 14776 27896 14804
rect 27890 14764 27896 14776
rect 27948 14764 27954 14816
rect 28074 14804 28080 14816
rect 28035 14776 28080 14804
rect 28074 14764 28080 14776
rect 28132 14764 28138 14816
rect 28166 14764 28172 14816
rect 28224 14804 28230 14816
rect 33318 14804 33324 14816
rect 28224 14776 33324 14804
rect 28224 14764 28230 14776
rect 33318 14764 33324 14776
rect 33376 14804 33382 14816
rect 34609 14807 34667 14813
rect 34609 14804 34621 14807
rect 33376 14776 34621 14804
rect 33376 14764 33382 14776
rect 34609 14773 34621 14776
rect 34655 14773 34667 14807
rect 43254 14804 43260 14816
rect 43215 14776 43260 14804
rect 34609 14767 34667 14773
rect 43254 14764 43260 14776
rect 43312 14764 43318 14816
rect 44085 14807 44143 14813
rect 44085 14773 44097 14807
rect 44131 14804 44143 14807
rect 44174 14804 44180 14816
rect 44131 14776 44180 14804
rect 44131 14773 44143 14776
rect 44085 14767 44143 14773
rect 44174 14764 44180 14776
rect 44232 14764 44238 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 2682 14600 2688 14612
rect 2643 14572 2688 14600
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 5132 14572 5181 14600
rect 5132 14560 5138 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 10778 14600 10784 14612
rect 9640 14572 10784 14600
rect 9640 14560 9646 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 15470 14600 15476 14612
rect 13320 14572 15476 14600
rect 13320 14560 13326 14572
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16022 14600 16028 14612
rect 15795 14572 16028 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 16393 14603 16451 14609
rect 16393 14569 16405 14603
rect 16439 14569 16451 14603
rect 16574 14600 16580 14612
rect 16535 14572 16580 14600
rect 16393 14563 16451 14569
rect 11606 14532 11612 14544
rect 2746 14504 11612 14532
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 2746 14464 2774 14504
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 16132 14532 16160 14560
rect 16408 14532 16436 14563
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 18138 14600 18144 14612
rect 18099 14572 18144 14600
rect 18138 14560 18144 14572
rect 18196 14560 18202 14612
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 25958 14600 25964 14612
rect 18380 14572 25964 14600
rect 18380 14560 18386 14572
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 26697 14603 26755 14609
rect 26697 14569 26709 14603
rect 26743 14600 26755 14603
rect 27430 14600 27436 14612
rect 26743 14572 27436 14600
rect 26743 14569 26755 14572
rect 26697 14563 26755 14569
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 27890 14560 27896 14612
rect 27948 14600 27954 14612
rect 31202 14600 31208 14612
rect 27948 14572 31208 14600
rect 27948 14560 27954 14572
rect 31202 14560 31208 14572
rect 31260 14600 31266 14612
rect 31386 14600 31392 14612
rect 31260 14572 31392 14600
rect 31260 14560 31266 14572
rect 31386 14560 31392 14572
rect 31444 14560 31450 14612
rect 31941 14603 31999 14609
rect 31941 14569 31953 14603
rect 31987 14600 31999 14603
rect 32398 14600 32404 14612
rect 31987 14572 32404 14600
rect 31987 14569 31999 14572
rect 31941 14563 31999 14569
rect 32398 14560 32404 14572
rect 32456 14560 32462 14612
rect 33689 14603 33747 14609
rect 33689 14569 33701 14603
rect 33735 14600 33747 14603
rect 34054 14600 34060 14612
rect 33735 14572 34060 14600
rect 33735 14569 33747 14572
rect 33689 14563 33747 14569
rect 34054 14560 34060 14572
rect 34112 14560 34118 14612
rect 35894 14560 35900 14612
rect 35952 14600 35958 14612
rect 36173 14603 36231 14609
rect 36173 14600 36185 14603
rect 35952 14572 36185 14600
rect 35952 14560 35958 14572
rect 36173 14569 36185 14572
rect 36219 14569 36231 14603
rect 37366 14600 37372 14612
rect 37327 14572 37372 14600
rect 36173 14563 36231 14569
rect 37366 14560 37372 14572
rect 37424 14560 37430 14612
rect 37458 14560 37464 14612
rect 37516 14600 37522 14612
rect 37516 14572 37561 14600
rect 37516 14560 37522 14572
rect 38654 14560 38660 14612
rect 38712 14600 38718 14612
rect 40129 14603 40187 14609
rect 40129 14600 40141 14603
rect 38712 14572 40141 14600
rect 38712 14560 38718 14572
rect 40129 14569 40141 14572
rect 40175 14569 40187 14603
rect 40129 14563 40187 14569
rect 43438 14560 43444 14612
rect 43496 14600 43502 14612
rect 43625 14603 43683 14609
rect 43625 14600 43637 14603
rect 43496 14572 43637 14600
rect 43496 14560 43502 14572
rect 43625 14569 43637 14572
rect 43671 14569 43683 14603
rect 43625 14563 43683 14569
rect 15672 14504 16436 14532
rect 16960 14504 27292 14532
rect 7650 14464 7656 14476
rect 1719 14436 2774 14464
rect 7484 14436 7656 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 2866 14396 2872 14408
rect 2827 14368 2872 14396
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 5350 14396 5356 14408
rect 5311 14368 5356 14396
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 6730 14396 6736 14408
rect 5675 14368 6736 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 7484 14405 7512 14436
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 12253 14467 12311 14473
rect 12253 14464 12265 14467
rect 10520 14436 12265 14464
rect 10520 14408 10548 14436
rect 12253 14433 12265 14436
rect 12299 14433 12311 14467
rect 12253 14427 12311 14433
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 14366 14464 14372 14476
rect 12759 14436 12940 14464
rect 14327 14436 14372 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 5537 14263 5595 14269
rect 5537 14229 5549 14263
rect 5583 14260 5595 14263
rect 5626 14260 5632 14272
rect 5583 14232 5632 14260
rect 5583 14229 5595 14232
rect 5537 14223 5595 14229
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 7576 14260 7604 14359
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 10502 14396 10508 14408
rect 7800 14368 7845 14396
rect 10463 14368 10508 14396
rect 7800 14356 7806 14368
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10778 14396 10784 14408
rect 10739 14368 10784 14396
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 11195 14368 12817 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 7653 14331 7711 14337
rect 7653 14297 7665 14331
rect 7699 14297 7711 14331
rect 8202 14328 8208 14340
rect 7653 14291 7711 14297
rect 7852 14300 8208 14328
rect 7524 14232 7604 14260
rect 7668 14260 7696 14291
rect 7852 14260 7880 14300
rect 8202 14288 8208 14300
rect 8260 14288 8266 14340
rect 9490 14288 9496 14340
rect 9548 14328 9554 14340
rect 11164 14328 11192 14359
rect 12912 14328 12940 14436
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 15672 14408 15700 14504
rect 14636 14399 14694 14405
rect 14636 14365 14648 14399
rect 14682 14396 14694 14399
rect 15010 14396 15016 14408
rect 14682 14368 15016 14396
rect 14682 14365 14694 14368
rect 14636 14359 14694 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 9548 14300 11192 14328
rect 11256 14300 12940 14328
rect 9548 14288 9554 14300
rect 7668 14232 7880 14260
rect 7929 14263 7987 14269
rect 7524 14220 7530 14232
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 9582 14260 9588 14272
rect 7975 14232 9588 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11256 14260 11284 14300
rect 16022 14288 16028 14340
rect 16080 14328 16086 14340
rect 16209 14331 16267 14337
rect 16209 14328 16221 14331
rect 16080 14300 16221 14328
rect 16080 14288 16086 14300
rect 16209 14297 16221 14300
rect 16255 14297 16267 14331
rect 16425 14331 16483 14337
rect 16425 14328 16437 14331
rect 16209 14291 16267 14297
rect 16408 14297 16437 14328
rect 16471 14328 16483 14331
rect 16960 14328 16988 14504
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18288 14436 18429 14464
rect 18288 14424 18294 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18509 14467 18567 14473
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 18555 14436 22017 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 22005 14433 22017 14436
rect 22051 14464 22063 14467
rect 23198 14464 23204 14476
rect 22051 14436 23204 14464
rect 22051 14433 22063 14436
rect 22005 14427 22063 14433
rect 23198 14424 23204 14436
rect 23256 14424 23262 14476
rect 25038 14424 25044 14476
rect 25096 14424 25102 14476
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 26510 14464 26516 14476
rect 25271 14436 26516 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 27264 14464 27292 14504
rect 28258 14492 28264 14544
rect 28316 14532 28322 14544
rect 31662 14532 31668 14544
rect 28316 14504 31668 14532
rect 28316 14492 28322 14504
rect 31662 14492 31668 14504
rect 31720 14492 31726 14544
rect 39114 14532 39120 14544
rect 33980 14504 39120 14532
rect 27264 14436 27384 14464
rect 18322 14396 18328 14408
rect 18283 14368 18328 14396
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 18598 14396 18604 14408
rect 18559 14368 18604 14396
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 21358 14356 21364 14408
rect 21416 14396 21422 14408
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21416 14368 21649 14396
rect 21416 14356 21422 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 21729 14399 21787 14405
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 22922 14396 22928 14408
rect 21775 14368 22928 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 23014 14356 23020 14408
rect 23072 14396 23078 14408
rect 25056 14396 25084 14424
rect 25866 14396 25872 14408
rect 23072 14368 25872 14396
rect 23072 14356 23078 14368
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 26602 14396 26608 14408
rect 26563 14368 26608 14396
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14365 26847 14399
rect 27246 14396 27252 14408
rect 27207 14368 27252 14396
rect 26789 14359 26847 14365
rect 16471 14300 16988 14328
rect 16471 14297 16483 14300
rect 16408 14291 16483 14297
rect 10836 14232 11284 14260
rect 11793 14263 11851 14269
rect 10836 14220 10842 14232
rect 11793 14229 11805 14263
rect 11839 14260 11851 14263
rect 11974 14260 11980 14272
rect 11839 14232 11980 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12437 14263 12495 14269
rect 12437 14229 12449 14263
rect 12483 14260 12495 14263
rect 16408 14260 16436 14291
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 22097 14331 22155 14337
rect 20312 14300 21588 14328
rect 20312 14288 20318 14300
rect 21450 14260 21456 14272
rect 12483 14232 16436 14260
rect 21411 14232 21456 14260
rect 12483 14229 12495 14232
rect 12437 14223 12495 14229
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 21560 14260 21588 14300
rect 22097 14297 22109 14331
rect 22143 14328 22155 14331
rect 22186 14328 22192 14340
rect 22143 14300 22192 14328
rect 22143 14297 22155 14300
rect 22097 14291 22155 14297
rect 22186 14288 22192 14300
rect 22244 14288 22250 14340
rect 25041 14331 25099 14337
rect 25041 14297 25053 14331
rect 25087 14297 25099 14331
rect 25041 14291 25099 14297
rect 25056 14260 25084 14291
rect 21560 14232 25084 14260
rect 26804 14260 26832 14359
rect 27246 14356 27252 14368
rect 27304 14356 27310 14408
rect 27356 14328 27384 14436
rect 30374 14424 30380 14476
rect 30432 14464 30438 14476
rect 30745 14467 30803 14473
rect 30745 14464 30757 14467
rect 30432 14436 30757 14464
rect 30432 14424 30438 14436
rect 30745 14433 30757 14436
rect 30791 14433 30803 14467
rect 31018 14464 31024 14476
rect 30979 14436 31024 14464
rect 30745 14427 30803 14433
rect 31018 14424 31024 14436
rect 31076 14424 31082 14476
rect 33980 14464 34008 14504
rect 39114 14492 39120 14504
rect 39172 14492 39178 14544
rect 43714 14532 43720 14544
rect 43675 14504 43720 14532
rect 43714 14492 43720 14504
rect 43772 14492 43778 14544
rect 31128 14436 34008 14464
rect 31128 14408 31156 14436
rect 34054 14424 34060 14476
rect 34112 14464 34118 14476
rect 34238 14464 34244 14476
rect 34112 14436 34244 14464
rect 34112 14424 34118 14436
rect 34238 14424 34244 14436
rect 34296 14424 34302 14476
rect 37918 14464 37924 14476
rect 37108 14436 37924 14464
rect 27516 14399 27574 14405
rect 27516 14365 27528 14399
rect 27562 14396 27574 14399
rect 28074 14396 28080 14408
rect 27562 14368 28080 14396
rect 27562 14365 27574 14368
rect 27516 14359 27574 14365
rect 28074 14356 28080 14368
rect 28132 14356 28138 14408
rect 30834 14396 30840 14408
rect 30795 14368 30840 14396
rect 30834 14356 30840 14368
rect 30892 14356 30898 14408
rect 30929 14399 30987 14405
rect 30929 14365 30941 14399
rect 30975 14396 30987 14399
rect 31110 14396 31116 14408
rect 30975 14368 31116 14396
rect 30975 14365 30987 14368
rect 30929 14359 30987 14365
rect 31110 14356 31116 14368
rect 31168 14356 31174 14408
rect 31386 14356 31392 14408
rect 31444 14396 31450 14408
rect 31573 14399 31631 14405
rect 31573 14396 31585 14399
rect 31444 14368 31585 14396
rect 31444 14356 31450 14368
rect 31573 14365 31585 14368
rect 31619 14365 31631 14399
rect 31573 14359 31631 14365
rect 31662 14356 31668 14408
rect 31720 14396 31726 14408
rect 31757 14399 31815 14405
rect 31757 14396 31769 14399
rect 31720 14368 31769 14396
rect 31720 14356 31726 14368
rect 31757 14365 31769 14368
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 33505 14399 33563 14405
rect 33505 14365 33517 14399
rect 33551 14396 33563 14399
rect 33594 14396 33600 14408
rect 33551 14368 33600 14396
rect 33551 14365 33563 14368
rect 33505 14359 33563 14365
rect 33594 14356 33600 14368
rect 33652 14356 33658 14408
rect 36081 14399 36139 14405
rect 36081 14365 36093 14399
rect 36127 14396 36139 14399
rect 36354 14396 36360 14408
rect 36127 14368 36360 14396
rect 36127 14365 36139 14368
rect 36081 14359 36139 14365
rect 36354 14356 36360 14368
rect 36412 14396 36418 14408
rect 36722 14396 36728 14408
rect 36412 14368 36728 14396
rect 36412 14356 36418 14368
rect 36722 14356 36728 14368
rect 36780 14356 36786 14408
rect 36998 14396 37004 14408
rect 36959 14368 37004 14396
rect 36998 14356 37004 14368
rect 37056 14356 37062 14408
rect 37108 14405 37136 14436
rect 37918 14424 37924 14436
rect 37976 14464 37982 14476
rect 38470 14464 38476 14476
rect 37976 14436 38476 14464
rect 37976 14424 37982 14436
rect 38470 14424 38476 14436
rect 38528 14464 38534 14476
rect 40313 14467 40371 14473
rect 40313 14464 40325 14467
rect 38528 14436 40325 14464
rect 38528 14424 38534 14436
rect 40313 14433 40325 14436
rect 40359 14433 40371 14467
rect 40313 14427 40371 14433
rect 43254 14424 43260 14476
rect 43312 14464 43318 14476
rect 43901 14467 43959 14473
rect 43901 14464 43913 14467
rect 43312 14436 43913 14464
rect 43312 14424 43318 14436
rect 43901 14433 43913 14436
rect 43947 14433 43959 14467
rect 43901 14427 43959 14433
rect 37093 14399 37151 14405
rect 37093 14365 37105 14399
rect 37139 14365 37151 14399
rect 37093 14359 37151 14365
rect 37461 14399 37519 14405
rect 37461 14365 37473 14399
rect 37507 14365 37519 14399
rect 37461 14359 37519 14365
rect 40037 14399 40095 14405
rect 40037 14365 40049 14399
rect 40083 14396 40095 14399
rect 40862 14396 40868 14408
rect 40083 14368 40868 14396
rect 40083 14365 40095 14368
rect 40037 14359 40095 14365
rect 28718 14328 28724 14340
rect 27356 14300 28724 14328
rect 28718 14288 28724 14300
rect 28776 14288 28782 14340
rect 28810 14288 28816 14340
rect 28868 14328 28874 14340
rect 32766 14328 32772 14340
rect 28868 14300 32772 14328
rect 28868 14288 28874 14300
rect 32766 14288 32772 14300
rect 32824 14288 32830 14340
rect 35802 14328 35808 14340
rect 33612 14300 35808 14328
rect 27062 14260 27068 14272
rect 26804 14232 27068 14260
rect 27062 14220 27068 14232
rect 27120 14260 27126 14272
rect 28258 14260 28264 14272
rect 27120 14232 28264 14260
rect 27120 14220 27126 14232
rect 28258 14220 28264 14232
rect 28316 14260 28322 14272
rect 28629 14263 28687 14269
rect 28629 14260 28641 14263
rect 28316 14232 28641 14260
rect 28316 14220 28322 14232
rect 28629 14229 28641 14232
rect 28675 14229 28687 14263
rect 28629 14223 28687 14229
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 30561 14263 30619 14269
rect 30561 14260 30573 14263
rect 30432 14232 30573 14260
rect 30432 14220 30438 14232
rect 30561 14229 30573 14232
rect 30607 14229 30619 14263
rect 30561 14223 30619 14229
rect 31018 14220 31024 14272
rect 31076 14260 31082 14272
rect 33612 14260 33640 14300
rect 35802 14288 35808 14300
rect 35860 14288 35866 14340
rect 37476 14328 37504 14359
rect 40862 14356 40868 14368
rect 40920 14356 40926 14408
rect 43625 14399 43683 14405
rect 43625 14365 43637 14399
rect 43671 14396 43683 14399
rect 44450 14396 44456 14408
rect 43671 14368 44456 14396
rect 43671 14365 43683 14368
rect 43625 14359 43683 14365
rect 44450 14356 44456 14368
rect 44508 14356 44514 14408
rect 46569 14399 46627 14405
rect 46569 14365 46581 14399
rect 46615 14396 46627 14399
rect 48406 14396 48412 14408
rect 46615 14368 48412 14396
rect 46615 14365 46627 14368
rect 46569 14359 46627 14365
rect 48406 14356 48412 14368
rect 48464 14396 48470 14408
rect 50157 14399 50215 14405
rect 50157 14396 50169 14399
rect 48464 14368 50169 14396
rect 48464 14356 48470 14368
rect 50157 14365 50169 14368
rect 50203 14365 50215 14399
rect 50157 14359 50215 14365
rect 53653 14399 53711 14405
rect 53653 14365 53665 14399
rect 53699 14365 53711 14399
rect 53653 14359 53711 14365
rect 53837 14399 53895 14405
rect 53837 14365 53849 14399
rect 53883 14396 53895 14399
rect 54018 14396 54024 14408
rect 53883 14368 54024 14396
rect 53883 14365 53895 14368
rect 53837 14359 53895 14365
rect 36096 14300 37504 14328
rect 31076 14232 33640 14260
rect 31076 14220 31082 14232
rect 33870 14220 33876 14272
rect 33928 14260 33934 14272
rect 36096 14260 36124 14300
rect 46290 14288 46296 14340
rect 46348 14328 46354 14340
rect 46814 14331 46872 14337
rect 46814 14328 46826 14331
rect 46348 14300 46826 14328
rect 46348 14288 46354 14300
rect 46814 14297 46826 14300
rect 46860 14297 46872 14331
rect 46814 14291 46872 14297
rect 50424 14331 50482 14337
rect 50424 14297 50436 14331
rect 50470 14328 50482 14331
rect 50614 14328 50620 14340
rect 50470 14300 50620 14328
rect 50470 14297 50482 14300
rect 50424 14291 50482 14297
rect 50614 14288 50620 14300
rect 50672 14288 50678 14340
rect 53668 14328 53696 14359
rect 54018 14356 54024 14368
rect 54076 14356 54082 14408
rect 54570 14328 54576 14340
rect 53668 14300 54576 14328
rect 54570 14288 54576 14300
rect 54628 14288 54634 14340
rect 33928 14232 36124 14260
rect 33928 14220 33934 14232
rect 36170 14220 36176 14272
rect 36228 14260 36234 14272
rect 36541 14263 36599 14269
rect 36541 14260 36553 14263
rect 36228 14232 36553 14260
rect 36228 14220 36234 14232
rect 36541 14229 36553 14232
rect 36587 14229 36599 14263
rect 36541 14223 36599 14229
rect 37185 14263 37243 14269
rect 37185 14229 37197 14263
rect 37231 14260 37243 14263
rect 37826 14260 37832 14272
rect 37231 14232 37832 14260
rect 37231 14229 37243 14232
rect 37185 14223 37243 14229
rect 37826 14220 37832 14232
rect 37884 14220 37890 14272
rect 40589 14263 40647 14269
rect 40589 14229 40601 14263
rect 40635 14260 40647 14263
rect 41046 14260 41052 14272
rect 40635 14232 41052 14260
rect 40635 14229 40647 14232
rect 40589 14223 40647 14229
rect 41046 14220 41052 14232
rect 41104 14220 41110 14272
rect 47946 14260 47952 14272
rect 47907 14232 47952 14260
rect 47946 14220 47952 14232
rect 48004 14220 48010 14272
rect 50154 14220 50160 14272
rect 50212 14260 50218 14272
rect 51537 14263 51595 14269
rect 51537 14260 51549 14263
rect 50212 14232 51549 14260
rect 50212 14220 50218 14232
rect 51537 14229 51549 14232
rect 51583 14229 51595 14263
rect 53742 14260 53748 14272
rect 53703 14232 53748 14260
rect 51537 14223 51595 14229
rect 53742 14220 53748 14232
rect 53800 14220 53806 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14056 2191 14059
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 2179 14028 3249 14056
rect 2179 14025 2191 14028
rect 2133 14019 2191 14025
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 12434 14056 12440 14068
rect 11011 14028 12440 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 14783 14059 14841 14065
rect 14783 14056 14795 14059
rect 13596 14028 14795 14056
rect 13596 14016 13602 14028
rect 14783 14025 14795 14028
rect 14829 14056 14841 14059
rect 15470 14056 15476 14068
rect 14829 14028 15476 14056
rect 14829 14025 14841 14028
rect 14783 14019 14841 14025
rect 15470 14016 15476 14028
rect 15528 14056 15534 14068
rect 15654 14056 15660 14068
rect 15528 14028 15660 14056
rect 15528 14016 15534 14028
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 23014 14056 23020 14068
rect 21416 14028 23020 14056
rect 21416 14016 21422 14028
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23198 14056 23204 14068
rect 23159 14028 23204 14056
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 24394 14016 24400 14068
rect 24452 14016 24458 14068
rect 24486 14016 24492 14068
rect 24544 14056 24550 14068
rect 28810 14056 28816 14068
rect 24544 14028 28816 14056
rect 24544 14016 24550 14028
rect 28810 14016 28816 14028
rect 28868 14016 28874 14068
rect 28920 14028 30604 14056
rect 6086 13988 6092 14000
rect 1412 13960 6092 13988
rect 1412 13929 1440 13960
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 10597 13991 10655 13997
rect 7800 13960 8432 13988
rect 7800 13948 7806 13960
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13889 1455 13923
rect 2314 13920 2320 13932
rect 2275 13892 2320 13920
rect 1397 13883 1455 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 5166 13920 5172 13932
rect 3191 13892 5172 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 7466 13880 7472 13932
rect 7524 13920 7530 13932
rect 7834 13920 7840 13932
rect 7524 13892 7840 13920
rect 7524 13880 7530 13892
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8202 13920 8208 13932
rect 8163 13892 8208 13920
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 8404 13929 8432 13960
rect 10597 13957 10609 13991
rect 10643 13988 10655 13991
rect 11514 13988 11520 14000
rect 10643 13960 11520 13988
rect 10643 13957 10655 13960
rect 10597 13951 10655 13957
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 11606 13948 11612 14000
rect 11664 13988 11670 14000
rect 16298 13988 16304 14000
rect 11664 13960 16304 13988
rect 11664 13948 11670 13960
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 21450 13948 21456 14000
rect 21508 13988 21514 14000
rect 22066 13991 22124 13997
rect 22066 13988 22078 13991
rect 21508 13960 22078 13988
rect 21508 13948 21514 13960
rect 22066 13957 22078 13960
rect 22112 13957 22124 13991
rect 24412 13988 24440 14016
rect 24642 13991 24700 13997
rect 24642 13988 24654 13991
rect 24412 13960 24654 13988
rect 22066 13951 22124 13957
rect 24642 13957 24654 13960
rect 24688 13957 24700 13991
rect 27982 13988 27988 14000
rect 27895 13960 27988 13988
rect 24642 13951 24700 13957
rect 27982 13948 27988 13960
rect 28040 13988 28046 14000
rect 28920 13988 28948 14028
rect 28040 13960 28948 13988
rect 28040 13948 28046 13960
rect 30374 13948 30380 14000
rect 30432 13997 30438 14000
rect 30432 13991 30496 13997
rect 30432 13957 30450 13991
rect 30484 13957 30496 13991
rect 30576 13988 30604 14028
rect 30650 14016 30656 14068
rect 30708 14056 30714 14068
rect 31386 14056 31392 14068
rect 30708 14028 31392 14056
rect 30708 14016 30714 14028
rect 31386 14016 31392 14028
rect 31444 14056 31450 14068
rect 31573 14059 31631 14065
rect 31573 14056 31585 14059
rect 31444 14028 31585 14056
rect 31444 14016 31450 14028
rect 31573 14025 31585 14028
rect 31619 14025 31631 14059
rect 31573 14019 31631 14025
rect 32309 14059 32367 14065
rect 32309 14025 32321 14059
rect 32355 14056 32367 14059
rect 32766 14056 32772 14068
rect 32355 14028 32772 14056
rect 32355 14025 32367 14028
rect 32309 14019 32367 14025
rect 32766 14016 32772 14028
rect 32824 14016 32830 14068
rect 40221 14059 40279 14065
rect 40221 14025 40233 14059
rect 40267 14056 40279 14059
rect 46658 14056 46664 14068
rect 40267 14028 43852 14056
rect 46619 14028 46664 14056
rect 40267 14025 40279 14028
rect 40221 14019 40279 14025
rect 40129 13991 40187 13997
rect 40129 13988 40141 13991
rect 30576 13960 40141 13988
rect 30432 13951 30496 13957
rect 40129 13957 40141 13960
rect 40175 13988 40187 13991
rect 40310 13988 40316 14000
rect 40175 13960 40316 13988
rect 40175 13957 40187 13960
rect 40129 13951 40187 13957
rect 30432 13948 30438 13951
rect 40310 13948 40316 13960
rect 40368 13948 40374 14000
rect 40402 13948 40408 14000
rect 40460 13988 40466 14000
rect 40957 13991 41015 13997
rect 40957 13988 40969 13991
rect 40460 13960 40969 13988
rect 40460 13948 40466 13960
rect 40957 13957 40969 13960
rect 41003 13957 41015 13991
rect 40957 13951 41015 13957
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 3050 13812 3056 13864
rect 3108 13852 3114 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 3108 13824 3341 13852
rect 3108 13812 3114 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 8956 13852 8984 13883
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10560 13892 10793 13920
rect 10560 13880 10566 13892
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 11974 13920 11980 13932
rect 11935 13892 11980 13920
rect 10781 13883 10839 13889
rect 11974 13880 11980 13892
rect 12032 13920 12038 13932
rect 20254 13920 20260 13932
rect 12032 13892 20260 13920
rect 12032 13880 12038 13892
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 21821 13923 21879 13929
rect 21821 13889 21833 13923
rect 21867 13920 21879 13923
rect 21910 13920 21916 13932
rect 21867 13892 21916 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 21910 13880 21916 13892
rect 21968 13920 21974 13932
rect 23934 13920 23940 13932
rect 21968 13892 23940 13920
rect 21968 13880 21974 13892
rect 23934 13880 23940 13892
rect 23992 13920 23998 13932
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 23992 13892 24409 13920
rect 23992 13880 23998 13892
rect 24397 13889 24409 13892
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 27890 13920 27896 13932
rect 27847 13892 27896 13920
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 27890 13880 27896 13892
rect 27948 13880 27954 13932
rect 28718 13880 28724 13932
rect 28776 13920 28782 13932
rect 30282 13920 30288 13932
rect 28776 13892 30288 13920
rect 28776 13880 28782 13892
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 32122 13920 32128 13932
rect 32083 13892 32128 13920
rect 32122 13880 32128 13892
rect 32180 13880 32186 13932
rect 33686 13920 33692 13932
rect 33647 13892 33692 13920
rect 33686 13880 33692 13892
rect 33744 13880 33750 13932
rect 34057 13923 34115 13929
rect 34057 13889 34069 13923
rect 34103 13920 34115 13923
rect 34238 13920 34244 13932
rect 34103 13892 34244 13920
rect 34103 13889 34115 13892
rect 34057 13883 34115 13889
rect 34238 13880 34244 13892
rect 34296 13880 34302 13932
rect 34790 13929 34796 13932
rect 34784 13883 34796 13929
rect 34848 13920 34854 13932
rect 34848 13892 34884 13920
rect 34790 13880 34796 13883
rect 34848 13880 34854 13892
rect 35894 13880 35900 13932
rect 35952 13920 35958 13932
rect 36541 13923 36599 13929
rect 36541 13920 36553 13923
rect 35952 13892 36553 13920
rect 35952 13880 35958 13892
rect 36541 13889 36553 13892
rect 36587 13889 36599 13923
rect 36722 13920 36728 13932
rect 36683 13892 36728 13920
rect 36541 13883 36599 13889
rect 36722 13880 36728 13892
rect 36780 13880 36786 13932
rect 40773 13923 40831 13929
rect 40773 13920 40785 13923
rect 40696 13892 40785 13920
rect 7064 13824 8984 13852
rect 12253 13855 12311 13861
rect 7064 13812 7070 13824
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 13078 13852 13084 13864
rect 12299 13824 13084 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13504 13824 13553 13852
rect 13504 13812 13510 13824
rect 13541 13821 13553 13824
rect 13587 13852 13599 13855
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 13587 13824 14565 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 14553 13821 14565 13824
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 16206 13852 16212 13864
rect 15896 13824 16212 13852
rect 15896 13812 15902 13824
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 26326 13812 26332 13864
rect 26384 13852 26390 13864
rect 27246 13852 27252 13864
rect 26384 13824 27252 13852
rect 26384 13812 26390 13824
rect 27246 13812 27252 13824
rect 27304 13852 27310 13864
rect 29270 13852 29276 13864
rect 27304 13824 29276 13852
rect 27304 13812 27310 13824
rect 29270 13812 29276 13824
rect 29328 13852 29334 13864
rect 30190 13852 30196 13864
rect 29328 13824 30196 13852
rect 29328 13812 29334 13824
rect 30190 13812 30196 13824
rect 30248 13812 30254 13864
rect 34514 13812 34520 13864
rect 34572 13852 34578 13864
rect 36633 13855 36691 13861
rect 36633 13852 36645 13855
rect 34572 13824 34617 13852
rect 36556 13824 36645 13852
rect 34572 13812 34578 13824
rect 36556 13796 36584 13824
rect 36633 13821 36645 13824
rect 36679 13852 36691 13855
rect 38746 13852 38752 13864
rect 36679 13824 38752 13852
rect 36679 13821 36691 13824
rect 36633 13815 36691 13821
rect 38746 13812 38752 13824
rect 38804 13812 38810 13864
rect 40034 13812 40040 13864
rect 40092 13852 40098 13864
rect 40696 13852 40724 13892
rect 40773 13889 40785 13892
rect 40819 13889 40831 13923
rect 41046 13920 41052 13932
rect 41007 13892 41052 13920
rect 40773 13883 40831 13889
rect 41046 13880 41052 13892
rect 41104 13880 41110 13932
rect 43824 13920 43852 14028
rect 46658 14016 46664 14028
rect 46716 14016 46722 14068
rect 50614 14056 50620 14068
rect 50575 14028 50620 14056
rect 50614 14016 50620 14028
rect 50672 14016 50678 14068
rect 44450 13948 44456 14000
rect 44508 13988 44514 14000
rect 45465 13991 45523 13997
rect 44508 13960 45416 13988
rect 44508 13948 44514 13960
rect 45002 13920 45008 13932
rect 43824 13892 45008 13920
rect 45002 13880 45008 13892
rect 45060 13920 45066 13932
rect 45281 13923 45339 13929
rect 45281 13920 45293 13923
rect 45060 13892 45293 13920
rect 45060 13880 45066 13892
rect 45281 13889 45293 13892
rect 45327 13889 45339 13923
rect 45388 13920 45416 13960
rect 45465 13957 45477 13991
rect 45511 13988 45523 13991
rect 53190 13988 53196 14000
rect 45511 13960 53196 13988
rect 45511 13957 45523 13960
rect 45465 13951 45523 13957
rect 53190 13948 53196 13960
rect 53248 13948 53254 14000
rect 53460 13991 53518 13997
rect 53460 13957 53472 13991
rect 53506 13988 53518 13991
rect 53742 13988 53748 14000
rect 53506 13960 53748 13988
rect 53506 13957 53518 13960
rect 53460 13951 53518 13957
rect 53742 13948 53748 13960
rect 53800 13948 53806 14000
rect 46569 13923 46627 13929
rect 46569 13920 46581 13923
rect 45388 13892 46581 13920
rect 45281 13883 45339 13889
rect 46569 13889 46581 13892
rect 46615 13889 46627 13923
rect 50522 13920 50528 13932
rect 50483 13892 50528 13920
rect 46569 13883 46627 13889
rect 50522 13880 50528 13892
rect 50580 13880 50586 13932
rect 50614 13880 50620 13932
rect 50672 13920 50678 13932
rect 50709 13923 50767 13929
rect 50709 13920 50721 13923
rect 50672 13892 50721 13920
rect 50672 13880 50678 13892
rect 50709 13889 50721 13892
rect 50755 13889 50767 13923
rect 50709 13883 50767 13889
rect 41414 13852 41420 13864
rect 40092 13824 40724 13852
rect 40092 13812 40098 13824
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 17218 13784 17224 13796
rect 1912 13756 17224 13784
rect 1912 13744 1918 13756
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 21634 13784 21640 13796
rect 17368 13756 21640 13784
rect 17368 13744 17374 13756
rect 21634 13744 21640 13756
rect 21692 13744 21698 13796
rect 25866 13744 25872 13796
rect 25924 13784 25930 13796
rect 28994 13784 29000 13796
rect 25924 13756 29000 13784
rect 25924 13744 25930 13756
rect 28994 13744 29000 13756
rect 29052 13744 29058 13796
rect 36538 13744 36544 13796
rect 36596 13744 36602 13796
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 2777 13719 2835 13725
rect 2777 13685 2789 13719
rect 2823 13716 2835 13719
rect 3050 13716 3056 13728
rect 2823 13688 3056 13716
rect 2823 13685 2835 13688
rect 2777 13679 2835 13685
rect 3050 13676 3056 13688
rect 3108 13676 3114 13728
rect 9033 13719 9091 13725
rect 9033 13685 9045 13719
rect 9079 13716 9091 13719
rect 11698 13716 11704 13728
rect 9079 13688 11704 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 11698 13676 11704 13688
rect 11756 13716 11762 13728
rect 12342 13716 12348 13728
rect 11756 13688 12348 13716
rect 11756 13676 11762 13688
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 18138 13716 18144 13728
rect 13872 13688 18144 13716
rect 13872 13676 13878 13688
rect 18138 13676 18144 13688
rect 18196 13716 18202 13728
rect 19242 13716 19248 13728
rect 18196 13688 19248 13716
rect 18196 13676 18202 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 21818 13716 21824 13728
rect 20864 13688 21824 13716
rect 20864 13676 20870 13688
rect 21818 13676 21824 13688
rect 21876 13716 21882 13728
rect 25682 13716 25688 13728
rect 21876 13688 25688 13716
rect 21876 13676 21882 13688
rect 25682 13676 25688 13688
rect 25740 13676 25746 13728
rect 25777 13719 25835 13725
rect 25777 13685 25789 13719
rect 25823 13716 25835 13719
rect 26050 13716 26056 13728
rect 25823 13688 26056 13716
rect 25823 13685 25835 13688
rect 25777 13679 25835 13685
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 27982 13676 27988 13728
rect 28040 13716 28046 13728
rect 34238 13716 34244 13728
rect 28040 13688 34244 13716
rect 28040 13676 28046 13688
rect 34238 13676 34244 13688
rect 34296 13676 34302 13728
rect 35894 13716 35900 13728
rect 35855 13688 35900 13716
rect 35894 13676 35900 13688
rect 35952 13676 35958 13728
rect 40696 13716 40724 13824
rect 40788 13824 41420 13852
rect 40788 13793 40816 13824
rect 41414 13812 41420 13824
rect 41472 13812 41478 13864
rect 44358 13812 44364 13864
rect 44416 13852 44422 13864
rect 45097 13855 45155 13861
rect 45097 13852 45109 13855
rect 44416 13824 45109 13852
rect 44416 13812 44422 13824
rect 45097 13821 45109 13824
rect 45143 13821 45155 13855
rect 45097 13815 45155 13821
rect 46845 13855 46903 13861
rect 46845 13821 46857 13855
rect 46891 13852 46903 13855
rect 47946 13852 47952 13864
rect 46891 13824 47952 13852
rect 46891 13821 46903 13824
rect 46845 13815 46903 13821
rect 47946 13812 47952 13824
rect 48004 13812 48010 13864
rect 52638 13812 52644 13864
rect 52696 13852 52702 13864
rect 53098 13852 53104 13864
rect 52696 13824 53104 13852
rect 52696 13812 52702 13824
rect 53098 13812 53104 13824
rect 53156 13852 53162 13864
rect 53193 13855 53251 13861
rect 53193 13852 53205 13855
rect 53156 13824 53205 13852
rect 53156 13812 53162 13824
rect 53193 13821 53205 13824
rect 53239 13821 53251 13855
rect 53193 13815 53251 13821
rect 40773 13787 40831 13793
rect 40773 13753 40785 13787
rect 40819 13753 40831 13787
rect 40773 13747 40831 13753
rect 45462 13716 45468 13728
rect 40696 13688 45468 13716
rect 45462 13676 45468 13688
rect 45520 13676 45526 13728
rect 46198 13716 46204 13728
rect 46159 13688 46204 13716
rect 46198 13676 46204 13688
rect 46256 13676 46262 13728
rect 54110 13676 54116 13728
rect 54168 13716 54174 13728
rect 54573 13719 54631 13725
rect 54573 13716 54585 13719
rect 54168 13688 54585 13716
rect 54168 13676 54174 13688
rect 54573 13685 54585 13688
rect 54619 13685 54631 13719
rect 54573 13679 54631 13685
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 6917 13515 6975 13521
rect 6917 13481 6929 13515
rect 6963 13512 6975 13515
rect 7374 13512 7380 13524
rect 6963 13484 7380 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 11057 13515 11115 13521
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 12618 13512 12624 13524
rect 11103 13484 12624 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 17218 13472 17224 13524
rect 17276 13512 17282 13524
rect 22830 13512 22836 13524
rect 17276 13484 22836 13512
rect 17276 13472 17282 13484
rect 22830 13472 22836 13484
rect 22888 13472 22894 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 28169 13515 28227 13521
rect 28169 13512 28181 13515
rect 25740 13484 28181 13512
rect 25740 13472 25746 13484
rect 28169 13481 28181 13484
rect 28215 13481 28227 13515
rect 28169 13475 28227 13481
rect 28813 13515 28871 13521
rect 28813 13481 28825 13515
rect 28859 13512 28871 13515
rect 29914 13512 29920 13524
rect 28859 13484 29920 13512
rect 28859 13481 28871 13484
rect 28813 13475 28871 13481
rect 5166 13444 5172 13456
rect 5079 13416 5172 13444
rect 5166 13404 5172 13416
rect 5224 13444 5230 13456
rect 7926 13444 7932 13456
rect 5224 13416 7932 13444
rect 5224 13404 5230 13416
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 10321 13447 10379 13453
rect 10321 13444 10333 13447
rect 8628 13416 10333 13444
rect 8628 13404 8634 13416
rect 10321 13413 10333 13416
rect 10367 13444 10379 13447
rect 10502 13444 10508 13456
rect 10367 13416 10508 13444
rect 10367 13413 10379 13416
rect 10321 13407 10379 13413
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18693 13447 18751 13453
rect 18693 13444 18705 13447
rect 18564 13416 18705 13444
rect 18564 13404 18570 13416
rect 18693 13413 18705 13416
rect 18739 13413 18751 13447
rect 26786 13444 26792 13456
rect 18693 13407 18751 13413
rect 18800 13416 19334 13444
rect 3786 13376 3792 13388
rect 3747 13348 3792 13376
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7558 13376 7564 13388
rect 7423 13348 7564 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 9490 13336 9496 13388
rect 9548 13376 9554 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9548 13348 10057 13376
rect 9548 13336 9554 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 13262 13336 13268 13388
rect 13320 13376 13326 13388
rect 13320 13348 17448 13376
rect 13320 13336 13326 13348
rect 3050 13308 3056 13320
rect 3011 13280 3056 13308
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 7190 13308 7196 13320
rect 6595 13280 7196 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7650 13308 7656 13320
rect 7611 13280 7656 13308
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 2222 13240 2228 13252
rect 2183 13212 2228 13240
rect 2222 13200 2228 13212
rect 2280 13200 2286 13252
rect 4034 13243 4092 13249
rect 4034 13240 4046 13243
rect 2884 13212 4046 13240
rect 2884 13181 2912 13212
rect 4034 13209 4046 13212
rect 4080 13209 4092 13243
rect 4034 13203 4092 13209
rect 6733 13243 6791 13249
rect 6733 13209 6745 13243
rect 6779 13240 6791 13243
rect 7098 13240 7104 13252
rect 6779 13212 7104 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 7098 13200 7104 13212
rect 7156 13240 7162 13252
rect 7558 13240 7564 13252
rect 7156 13212 7564 13240
rect 7156 13200 7162 13212
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 2869 13175 2927 13181
rect 2869 13141 2881 13175
rect 2915 13141 2927 13175
rect 2869 13135 2927 13141
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9508 13172 9536 13336
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 14108 13317 14136 13348
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 9640 13280 10977 13308
rect 9640 13268 9646 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 17276 13280 17325 13308
rect 17276 13268 17282 13280
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17420 13308 17448 13348
rect 18800 13308 18828 13416
rect 17420 13280 18828 13308
rect 17313 13271 17371 13277
rect 17580 13243 17638 13249
rect 17580 13209 17592 13243
rect 17626 13240 17638 13243
rect 17954 13240 17960 13252
rect 17626 13212 17960 13240
rect 17626 13209 17638 13212
rect 17580 13203 17638 13209
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 19306 13240 19334 13416
rect 20548 13416 26792 13444
rect 20162 13336 20168 13388
rect 20220 13376 20226 13388
rect 20548 13385 20576 13416
rect 26786 13404 26792 13416
rect 26844 13404 26850 13456
rect 28184 13444 28212 13475
rect 29914 13472 29920 13484
rect 29972 13512 29978 13524
rect 30098 13512 30104 13524
rect 29972 13484 30104 13512
rect 29972 13472 29978 13484
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 30469 13515 30527 13521
rect 30469 13481 30481 13515
rect 30515 13512 30527 13515
rect 30834 13512 30840 13524
rect 30515 13484 30840 13512
rect 30515 13481 30527 13484
rect 30469 13475 30527 13481
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 32309 13515 32367 13521
rect 32309 13481 32321 13515
rect 32355 13512 32367 13515
rect 32858 13512 32864 13524
rect 32355 13484 32864 13512
rect 32355 13481 32367 13484
rect 32309 13475 32367 13481
rect 32858 13472 32864 13484
rect 32916 13472 32922 13524
rect 33410 13512 33416 13524
rect 33371 13484 33416 13512
rect 33410 13472 33416 13484
rect 33468 13472 33474 13524
rect 34790 13472 34796 13524
rect 34848 13512 34854 13524
rect 35069 13515 35127 13521
rect 35069 13512 35081 13515
rect 34848 13484 35081 13512
rect 34848 13472 34854 13484
rect 35069 13481 35081 13484
rect 35115 13481 35127 13515
rect 36354 13512 36360 13524
rect 36315 13484 36360 13512
rect 35069 13475 35127 13481
rect 36354 13472 36360 13484
rect 36412 13472 36418 13524
rect 36633 13515 36691 13521
rect 36633 13481 36645 13515
rect 36679 13512 36691 13515
rect 36722 13512 36728 13524
rect 36679 13484 36728 13512
rect 36679 13481 36691 13484
rect 36633 13475 36691 13481
rect 36722 13472 36728 13484
rect 36780 13512 36786 13524
rect 36998 13512 37004 13524
rect 36780 13484 37004 13512
rect 36780 13472 36786 13484
rect 36998 13472 37004 13484
rect 37056 13472 37062 13524
rect 40221 13515 40279 13521
rect 40221 13481 40233 13515
rect 40267 13512 40279 13515
rect 44082 13512 44088 13524
rect 40267 13484 41000 13512
rect 44043 13484 44088 13512
rect 40267 13481 40279 13484
rect 40221 13475 40279 13481
rect 32122 13444 32128 13456
rect 28184 13416 32128 13444
rect 32122 13404 32128 13416
rect 32180 13404 32186 13456
rect 34238 13404 34244 13456
rect 34296 13444 34302 13456
rect 36814 13444 36820 13456
rect 34296 13416 36820 13444
rect 34296 13404 34302 13416
rect 36814 13404 36820 13416
rect 36872 13404 36878 13456
rect 20533 13379 20591 13385
rect 20533 13376 20545 13379
rect 20220 13348 20545 13376
rect 20220 13336 20226 13348
rect 20533 13345 20545 13348
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 21726 13336 21732 13388
rect 21784 13376 21790 13388
rect 21784 13348 22600 13376
rect 21784 13336 21790 13348
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19484 13280 19809 13308
rect 19484 13268 19490 13280
rect 19797 13277 19809 13280
rect 19843 13308 19855 13311
rect 20070 13308 20076 13320
rect 19843 13280 20076 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20254 13308 20260 13320
rect 20215 13280 20260 13308
rect 20254 13268 20260 13280
rect 20312 13308 20318 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 20312 13280 21281 13308
rect 20312 13268 20318 13280
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 21450 13268 21456 13320
rect 21508 13308 21514 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21508 13280 21557 13308
rect 21508 13268 21514 13280
rect 21545 13277 21557 13280
rect 21591 13308 21603 13311
rect 22094 13308 22100 13320
rect 21591 13280 22100 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22572 13317 22600 13348
rect 28092 13348 28948 13376
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 22557 13271 22615 13277
rect 22741 13311 22799 13317
rect 22741 13277 22753 13311
rect 22787 13308 22799 13311
rect 22830 13308 22836 13320
rect 22787 13280 22836 13308
rect 22787 13277 22799 13280
rect 22741 13271 22799 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13308 24639 13311
rect 24670 13308 24676 13320
rect 24627 13280 24676 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 24854 13308 24860 13320
rect 24815 13280 24860 13308
rect 24854 13268 24860 13280
rect 24912 13268 24918 13320
rect 25041 13311 25099 13317
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 26602 13308 26608 13320
rect 25087 13280 26608 13308
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 27890 13240 27896 13252
rect 19306 13212 27896 13240
rect 27890 13200 27896 13212
rect 27948 13240 27954 13252
rect 28092 13249 28120 13348
rect 28718 13308 28724 13320
rect 28679 13280 28724 13308
rect 28718 13268 28724 13280
rect 28776 13268 28782 13320
rect 28920 13317 28948 13348
rect 28994 13336 29000 13388
rect 29052 13376 29058 13388
rect 34790 13376 34796 13388
rect 29052 13348 34796 13376
rect 29052 13336 29058 13348
rect 34790 13336 34796 13348
rect 34848 13376 34854 13388
rect 34848 13348 35296 13376
rect 34848 13336 34854 13348
rect 28905 13311 28963 13317
rect 28905 13277 28917 13311
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 29362 13268 29368 13320
rect 29420 13308 29426 13320
rect 30650 13308 30656 13320
rect 29420 13280 30656 13308
rect 29420 13268 29426 13280
rect 30650 13268 30656 13280
rect 30708 13268 30714 13320
rect 30926 13308 30932 13320
rect 30887 13280 30932 13308
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 32122 13308 32128 13320
rect 32083 13280 32128 13308
rect 32122 13268 32128 13280
rect 32180 13268 32186 13320
rect 35268 13317 35296 13348
rect 35253 13311 35311 13317
rect 35253 13277 35265 13311
rect 35299 13277 35311 13311
rect 35253 13271 35311 13277
rect 35529 13311 35587 13317
rect 35529 13277 35541 13311
rect 35575 13308 35587 13311
rect 36078 13308 36084 13320
rect 35575 13280 36084 13308
rect 35575 13277 35587 13280
rect 35529 13271 35587 13277
rect 36078 13268 36084 13280
rect 36136 13268 36142 13320
rect 36173 13311 36231 13317
rect 36173 13277 36185 13311
rect 36219 13277 36231 13311
rect 36173 13271 36231 13277
rect 28077 13243 28135 13249
rect 28077 13240 28089 13243
rect 27948 13212 28089 13240
rect 27948 13200 27954 13212
rect 28077 13209 28089 13212
rect 28123 13209 28135 13243
rect 28077 13203 28135 13209
rect 28166 13200 28172 13252
rect 28224 13240 28230 13252
rect 33134 13240 33140 13252
rect 28224 13212 33140 13240
rect 28224 13200 28230 13212
rect 33134 13200 33140 13212
rect 33192 13200 33198 13252
rect 35437 13243 35495 13249
rect 35437 13209 35449 13243
rect 35483 13240 35495 13243
rect 35894 13240 35900 13252
rect 35483 13212 35900 13240
rect 35483 13209 35495 13212
rect 35437 13203 35495 13209
rect 35894 13200 35900 13212
rect 35952 13240 35958 13252
rect 36188 13240 36216 13271
rect 36262 13268 36268 13320
rect 36320 13308 36326 13320
rect 36906 13308 36912 13320
rect 36320 13280 36912 13308
rect 36320 13268 36326 13280
rect 36906 13268 36912 13280
rect 36964 13268 36970 13320
rect 39758 13268 39764 13320
rect 39816 13308 39822 13320
rect 39945 13311 40003 13317
rect 39945 13308 39957 13311
rect 39816 13280 39957 13308
rect 39816 13268 39822 13280
rect 39945 13277 39957 13280
rect 39991 13308 40003 13311
rect 40678 13308 40684 13320
rect 39991 13280 40684 13308
rect 39991 13277 40003 13280
rect 39945 13271 40003 13277
rect 40678 13268 40684 13280
rect 40736 13268 40742 13320
rect 35952 13212 36216 13240
rect 35952 13200 35958 13212
rect 40972 13184 41000 13484
rect 44082 13472 44088 13484
rect 44140 13472 44146 13524
rect 44450 13512 44456 13524
rect 44411 13484 44456 13512
rect 44450 13472 44456 13484
rect 44508 13472 44514 13524
rect 46201 13515 46259 13521
rect 46201 13481 46213 13515
rect 46247 13512 46259 13515
rect 46290 13512 46296 13524
rect 46247 13484 46296 13512
rect 46247 13481 46259 13484
rect 46201 13475 46259 13481
rect 46290 13472 46296 13484
rect 46348 13472 46354 13524
rect 50433 13515 50491 13521
rect 50433 13481 50445 13515
rect 50479 13512 50491 13515
rect 50522 13512 50528 13524
rect 50479 13484 50528 13512
rect 50479 13481 50491 13484
rect 50433 13475 50491 13481
rect 50522 13472 50528 13484
rect 50580 13472 50586 13524
rect 54570 13512 54576 13524
rect 54531 13484 54576 13512
rect 54570 13472 54576 13484
rect 54628 13472 54634 13524
rect 45462 13404 45468 13456
rect 45520 13444 45526 13456
rect 45520 13416 46428 13444
rect 45520 13404 45526 13416
rect 41138 13376 41144 13388
rect 41099 13348 41144 13376
rect 41138 13336 41144 13348
rect 41196 13336 41202 13388
rect 44174 13376 44180 13388
rect 44135 13348 44180 13376
rect 44174 13336 44180 13348
rect 44232 13336 44238 13388
rect 41414 13317 41420 13320
rect 41408 13308 41420 13317
rect 41375 13280 41420 13308
rect 41408 13271 41420 13280
rect 41414 13268 41420 13271
rect 41472 13268 41478 13320
rect 44269 13311 44327 13317
rect 44269 13277 44281 13311
rect 44315 13308 44327 13311
rect 44358 13308 44364 13320
rect 44315 13280 44364 13308
rect 44315 13277 44327 13280
rect 44269 13271 44327 13277
rect 44358 13268 44364 13280
rect 44416 13268 44422 13320
rect 46198 13308 46204 13320
rect 46159 13280 46204 13308
rect 46198 13268 46204 13280
rect 46256 13268 46262 13320
rect 46400 13317 46428 13416
rect 48038 13404 48044 13456
rect 48096 13444 48102 13456
rect 48096 13416 54708 13444
rect 48096 13404 48102 13416
rect 50540 13385 50568 13416
rect 54680 13385 54708 13416
rect 50525 13379 50583 13385
rect 49344 13348 50384 13376
rect 46385 13311 46443 13317
rect 46385 13277 46397 13311
rect 46431 13277 46443 13311
rect 49142 13308 49148 13320
rect 49103 13280 49148 13308
rect 46385 13271 46443 13277
rect 49142 13268 49148 13280
rect 49200 13268 49206 13320
rect 49344 13317 49372 13348
rect 49329 13311 49387 13317
rect 49329 13277 49341 13311
rect 49375 13277 49387 13311
rect 49329 13271 49387 13277
rect 50154 13268 50160 13320
rect 50212 13308 50218 13320
rect 50356 13317 50384 13348
rect 50525 13345 50537 13379
rect 50571 13345 50583 13379
rect 54481 13379 54539 13385
rect 54481 13376 54493 13379
rect 50525 13339 50583 13345
rect 53760 13348 54493 13376
rect 53760 13320 53788 13348
rect 54481 13345 54493 13348
rect 54527 13345 54539 13379
rect 54481 13339 54539 13345
rect 54665 13379 54723 13385
rect 54665 13345 54677 13379
rect 54711 13376 54723 13379
rect 54938 13376 54944 13388
rect 54711 13348 54944 13376
rect 54711 13345 54723 13348
rect 54665 13339 54723 13345
rect 54938 13336 54944 13348
rect 54996 13336 55002 13388
rect 50249 13311 50307 13317
rect 50249 13308 50261 13311
rect 50212 13280 50261 13308
rect 50212 13268 50218 13280
rect 50249 13277 50261 13280
rect 50295 13277 50307 13311
rect 50249 13271 50307 13277
rect 50341 13311 50399 13317
rect 50341 13277 50353 13311
rect 50387 13308 50399 13311
rect 50982 13308 50988 13320
rect 50387 13280 50988 13308
rect 50387 13277 50399 13280
rect 50341 13271 50399 13277
rect 50982 13268 50988 13280
rect 51040 13268 51046 13320
rect 53653 13311 53711 13317
rect 53653 13277 53665 13311
rect 53699 13277 53711 13311
rect 53653 13271 53711 13277
rect 43809 13243 43867 13249
rect 43809 13240 43821 13243
rect 42536 13212 43821 13240
rect 10502 13172 10508 13184
rect 9456 13144 9536 13172
rect 10463 13144 10508 13172
rect 9456 13132 9462 13144
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 13964 13144 14289 13172
rect 13964 13132 13970 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14277 13135 14335 13141
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 18690 13172 18696 13184
rect 16172 13144 18696 13172
rect 16172 13132 16178 13144
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 22741 13175 22799 13181
rect 22741 13141 22753 13175
rect 22787 13172 22799 13175
rect 22922 13172 22928 13184
rect 22787 13144 22928 13172
rect 22787 13141 22799 13144
rect 22741 13135 22799 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 24394 13132 24400 13184
rect 24452 13172 24458 13184
rect 24765 13175 24823 13181
rect 24765 13172 24777 13175
rect 24452 13144 24777 13172
rect 24452 13132 24458 13144
rect 24765 13141 24777 13144
rect 24811 13141 24823 13175
rect 24765 13135 24823 13141
rect 26510 13132 26516 13184
rect 26568 13172 26574 13184
rect 28350 13172 28356 13184
rect 26568 13144 28356 13172
rect 26568 13132 26574 13144
rect 28350 13132 28356 13144
rect 28408 13172 28414 13184
rect 28902 13172 28908 13184
rect 28408 13144 28908 13172
rect 28408 13132 28414 13144
rect 28902 13132 28908 13144
rect 28960 13172 28966 13184
rect 29270 13172 29276 13184
rect 28960 13144 29276 13172
rect 28960 13132 28966 13144
rect 29270 13132 29276 13144
rect 29328 13132 29334 13184
rect 30837 13175 30895 13181
rect 30837 13141 30849 13175
rect 30883 13172 30895 13175
rect 31662 13172 31668 13184
rect 30883 13144 31668 13172
rect 30883 13141 30895 13144
rect 30837 13135 30895 13141
rect 31662 13132 31668 13144
rect 31720 13132 31726 13184
rect 40402 13172 40408 13184
rect 40363 13144 40408 13172
rect 40402 13132 40408 13144
rect 40460 13132 40466 13184
rect 40954 13132 40960 13184
rect 41012 13172 41018 13184
rect 42536 13181 42564 13212
rect 43809 13209 43821 13212
rect 43855 13240 43867 13243
rect 44634 13240 44640 13252
rect 43855 13212 44640 13240
rect 43855 13209 43867 13212
rect 43809 13203 43867 13209
rect 44634 13200 44640 13212
rect 44692 13200 44698 13252
rect 53668 13240 53696 13271
rect 53742 13268 53748 13320
rect 53800 13308 53806 13320
rect 54389 13311 54447 13317
rect 53800 13280 53845 13308
rect 53800 13268 53806 13280
rect 54389 13277 54401 13311
rect 54435 13277 54447 13311
rect 54389 13271 54447 13277
rect 54110 13240 54116 13252
rect 53668 13212 54116 13240
rect 54110 13200 54116 13212
rect 54168 13240 54174 13252
rect 54404 13240 54432 13271
rect 54168 13212 54432 13240
rect 54168 13200 54174 13212
rect 42521 13175 42579 13181
rect 42521 13172 42533 13175
rect 41012 13144 42533 13172
rect 41012 13132 41018 13144
rect 42521 13141 42533 13144
rect 42567 13141 42579 13175
rect 49234 13172 49240 13184
rect 49195 13144 49240 13172
rect 42521 13135 42579 13141
rect 49234 13132 49240 13144
rect 49292 13132 49298 13184
rect 53929 13175 53987 13181
rect 53929 13141 53941 13175
rect 53975 13172 53987 13175
rect 54018 13172 54024 13184
rect 53975 13144 54024 13172
rect 53975 13141 53987 13144
rect 53929 13135 53987 13141
rect 54018 13132 54024 13144
rect 54076 13132 54082 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 7742 12968 7748 12980
rect 7239 12940 7748 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 9950 12968 9956 12980
rect 7800 12940 9812 12968
rect 9911 12940 9956 12968
rect 7800 12928 7806 12940
rect 5902 12860 5908 12912
rect 5960 12900 5966 12912
rect 9784 12900 9812 12940
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 17954 12968 17960 12980
rect 11716 12940 16252 12968
rect 17915 12940 17960 12968
rect 5960 12872 8524 12900
rect 9784 12872 10088 12900
rect 5960 12860 5966 12872
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 2682 12832 2688 12844
rect 2643 12804 2688 12832
rect 1397 12795 1455 12801
rect 1412 12764 1440 12795
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3326 12832 3332 12844
rect 3287 12804 3332 12832
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 7190 12832 7196 12844
rect 7151 12804 7196 12832
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7616 12804 7849 12832
rect 7616 12792 7622 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 3970 12764 3976 12776
rect 1412 12736 3976 12764
rect 3970 12724 3976 12736
rect 4028 12724 4034 12776
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7800 12736 8309 12764
rect 7800 12724 7806 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8496 12764 8524 12872
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 10060 12841 10088 12872
rect 9861 12835 9919 12841
rect 8628 12804 8673 12832
rect 8628 12792 8634 12804
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10502 12832 10508 12844
rect 10463 12804 10508 12832
rect 10045 12795 10103 12801
rect 9882 12764 9910 12795
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 10686 12832 10692 12844
rect 10647 12804 10692 12832
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11716 12841 11744 12940
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 13265 12903 13323 12909
rect 13265 12900 13277 12903
rect 12584 12872 13277 12900
rect 12584 12860 12590 12872
rect 13265 12869 13277 12872
rect 13311 12869 13323 12903
rect 15286 12900 15292 12912
rect 15247 12872 15292 12900
rect 13265 12863 13323 12869
rect 15286 12860 15292 12872
rect 15344 12860 15350 12912
rect 15505 12903 15563 12909
rect 15505 12900 15517 12903
rect 15488 12869 15517 12900
rect 15551 12900 15563 12903
rect 16114 12900 16120 12912
rect 15551 12872 16120 12900
rect 15551 12869 15563 12872
rect 15488 12863 15563 12869
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 10928 12804 11713 12832
rect 10928 12792 10934 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 11701 12795 11759 12801
rect 11808 12804 12449 12832
rect 10134 12764 10140 12776
rect 8496 12736 9812 12764
rect 9882 12736 10140 12764
rect 8297 12727 8355 12733
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 9784 12696 9812 12736
rect 10134 12724 10140 12736
rect 10192 12764 10198 12776
rect 10520 12764 10548 12792
rect 10192 12736 10548 12764
rect 10192 12724 10198 12736
rect 11808 12705 11836 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13357 12835 13415 12841
rect 13357 12832 13369 12835
rect 13136 12804 13369 12832
rect 13136 12792 13142 12804
rect 13357 12801 13369 12804
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 15013 12835 15071 12841
rect 15013 12801 15025 12835
rect 15059 12832 15071 12835
rect 15488 12832 15516 12863
rect 16114 12860 16120 12872
rect 16172 12860 16178 12912
rect 16224 12900 16252 12940
rect 17954 12928 17960 12940
rect 18012 12928 18018 12980
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 18506 12968 18512 12980
rect 18371 12940 18512 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 20993 12971 21051 12977
rect 18748 12940 20944 12968
rect 18748 12928 18754 12940
rect 19426 12900 19432 12912
rect 16224 12872 19432 12900
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 19978 12900 19984 12912
rect 19939 12872 19984 12900
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 20806 12900 20812 12912
rect 20767 12872 20812 12900
rect 20806 12860 20812 12872
rect 20864 12860 20870 12912
rect 20916 12900 20944 12940
rect 20993 12937 21005 12971
rect 21039 12968 21051 12971
rect 21450 12968 21456 12980
rect 21039 12940 21456 12968
rect 21039 12937 21051 12940
rect 20993 12931 21051 12937
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 24397 12971 24455 12977
rect 24397 12937 24409 12971
rect 24443 12968 24455 12971
rect 24854 12968 24860 12980
rect 24443 12940 24860 12968
rect 24443 12937 24455 12940
rect 24397 12931 24455 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 28184 12940 29224 12968
rect 27982 12900 27988 12912
rect 20916 12872 27988 12900
rect 27982 12860 27988 12872
rect 28040 12860 28046 12912
rect 28184 12900 28212 12940
rect 28350 12900 28356 12912
rect 28092 12872 28212 12900
rect 28311 12872 28356 12900
rect 28092 12844 28120 12872
rect 28350 12860 28356 12872
rect 28408 12860 28414 12912
rect 15059 12804 15516 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 18138 12792 18144 12844
rect 18196 12841 18202 12844
rect 18196 12835 18218 12841
rect 18206 12801 18218 12835
rect 18196 12795 18218 12801
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 19150 12832 19156 12844
rect 18463 12804 19156 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 18196 12792 18202 12795
rect 19150 12792 19156 12804
rect 19208 12832 19214 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19208 12804 20177 12832
rect 19208 12792 19214 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12832 24179 12835
rect 26050 12832 26056 12844
rect 24167 12804 26056 12832
rect 24167 12801 24179 12804
rect 24121 12795 24179 12801
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 28074 12832 28080 12844
rect 27987 12804 28080 12832
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 28258 12841 28264 12844
rect 28225 12835 28264 12841
rect 28225 12801 28237 12835
rect 28225 12795 28264 12801
rect 28258 12792 28264 12795
rect 28316 12792 28322 12844
rect 28442 12832 28448 12844
rect 28403 12804 28448 12832
rect 28442 12792 28448 12804
rect 28500 12792 28506 12844
rect 28583 12835 28641 12841
rect 28583 12801 28595 12835
rect 28629 12832 28641 12835
rect 28718 12832 28724 12844
rect 28629 12804 28724 12832
rect 28629 12801 28641 12804
rect 28583 12795 28641 12801
rect 28718 12792 28724 12804
rect 28776 12832 28782 12844
rect 29196 12841 29224 12940
rect 29270 12928 29276 12980
rect 29328 12928 29334 12980
rect 33134 12928 33140 12980
rect 33192 12968 33198 12980
rect 48038 12968 48044 12980
rect 33192 12940 48044 12968
rect 33192 12928 33198 12940
rect 48038 12928 48044 12940
rect 48096 12928 48102 12980
rect 50982 12968 50988 12980
rect 50943 12940 50988 12968
rect 50982 12928 50988 12940
rect 51040 12928 51046 12980
rect 52638 12928 52644 12980
rect 52696 12968 52702 12980
rect 55858 12968 55864 12980
rect 52696 12940 55864 12968
rect 52696 12928 52702 12940
rect 55858 12928 55864 12940
rect 55916 12928 55922 12980
rect 57241 12971 57299 12977
rect 57241 12937 57253 12971
rect 57287 12937 57299 12971
rect 57241 12931 57299 12937
rect 29288 12900 29316 12928
rect 29457 12903 29515 12909
rect 29457 12900 29469 12903
rect 29288 12872 29469 12900
rect 29457 12869 29469 12872
rect 29503 12869 29515 12903
rect 29457 12863 29515 12869
rect 29549 12903 29607 12909
rect 29549 12869 29561 12903
rect 29595 12900 29607 12903
rect 30098 12900 30104 12912
rect 29595 12872 30104 12900
rect 29595 12869 29607 12872
rect 29549 12863 29607 12869
rect 30098 12860 30104 12872
rect 30156 12860 30162 12912
rect 38565 12903 38623 12909
rect 38565 12869 38577 12903
rect 38611 12900 38623 12903
rect 40402 12900 40408 12912
rect 38611 12872 40408 12900
rect 38611 12869 38623 12872
rect 38565 12863 38623 12869
rect 40402 12860 40408 12872
rect 40460 12860 40466 12912
rect 44634 12900 44640 12912
rect 44595 12872 44640 12900
rect 44634 12860 44640 12872
rect 44692 12860 44698 12912
rect 47854 12860 47860 12912
rect 47912 12900 47918 12912
rect 47949 12903 48007 12909
rect 47949 12900 47961 12903
rect 47912 12872 47961 12900
rect 47912 12860 47918 12872
rect 47949 12869 47961 12872
rect 47995 12900 48007 12903
rect 48222 12900 48228 12912
rect 47995 12872 48228 12900
rect 47995 12869 48007 12872
rect 47949 12863 48007 12869
rect 48222 12860 48228 12872
rect 48280 12860 48286 12912
rect 49044 12903 49102 12909
rect 49044 12869 49056 12903
rect 49090 12900 49102 12903
rect 49234 12900 49240 12912
rect 49090 12872 49240 12900
rect 49090 12869 49102 12872
rect 49044 12863 49102 12869
rect 49234 12860 49240 12872
rect 49292 12860 49298 12912
rect 55490 12900 55496 12912
rect 53852 12872 55496 12900
rect 53852 12844 53880 12872
rect 29362 12841 29368 12844
rect 29181 12835 29239 12841
rect 28776 12804 28994 12832
rect 28776 12792 28782 12804
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12764 12679 12767
rect 13262 12764 13268 12776
rect 12667 12736 13268 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 19242 12724 19248 12776
rect 19300 12764 19306 12776
rect 24394 12764 24400 12776
rect 19300 12736 22094 12764
rect 24355 12736 24400 12764
rect 19300 12724 19306 12736
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 3191 12668 9674 12696
rect 9784 12668 11805 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 9646 12640 9674 12668
rect 11793 12665 11805 12668
rect 11839 12665 11851 12699
rect 11793 12659 11851 12665
rect 13081 12699 13139 12705
rect 13081 12665 13093 12699
rect 13127 12696 13139 12699
rect 13446 12696 13452 12708
rect 13127 12668 13452 12696
rect 13127 12665 13139 12668
rect 13081 12659 13139 12665
rect 13446 12656 13452 12668
rect 13504 12656 13510 12708
rect 14366 12656 14372 12708
rect 14424 12696 14430 12708
rect 14424 12668 16252 12696
rect 14424 12656 14430 12668
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2866 12628 2872 12640
rect 2547 12600 2872 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 9646 12600 9680 12640
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 10873 12631 10931 12637
rect 10873 12597 10885 12631
rect 10919 12628 10931 12631
rect 10962 12628 10968 12640
rect 10919 12600 10968 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13630 12628 13636 12640
rect 13587 12600 13636 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15654 12628 15660 12640
rect 15615 12600 15660 12628
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 16224 12628 16252 12668
rect 16298 12656 16304 12708
rect 16356 12696 16362 12708
rect 20441 12699 20499 12705
rect 20441 12696 20453 12699
rect 16356 12668 20453 12696
rect 16356 12656 16362 12668
rect 20441 12665 20453 12668
rect 20487 12696 20499 12699
rect 22066 12696 22094 12736
rect 24394 12724 24400 12736
rect 24452 12724 24458 12776
rect 28966 12764 28994 12804
rect 29181 12801 29193 12835
rect 29227 12801 29239 12835
rect 29181 12795 29239 12801
rect 29329 12835 29368 12841
rect 29329 12801 29341 12835
rect 29329 12795 29368 12801
rect 29362 12792 29368 12795
rect 29420 12792 29426 12844
rect 29646 12835 29704 12841
rect 29646 12832 29658 12835
rect 29472 12804 29658 12832
rect 29472 12764 29500 12804
rect 29646 12801 29658 12804
rect 29692 12801 29704 12835
rect 38746 12832 38752 12844
rect 38707 12804 38752 12832
rect 29646 12795 29704 12801
rect 38746 12792 38752 12804
rect 38804 12792 38810 12844
rect 39758 12832 39764 12844
rect 39719 12804 39764 12832
rect 39758 12792 39764 12804
rect 39816 12792 39822 12844
rect 39945 12835 40003 12841
rect 39945 12801 39957 12835
rect 39991 12832 40003 12835
rect 40954 12832 40960 12844
rect 39991 12804 40960 12832
rect 39991 12801 40003 12804
rect 39945 12795 40003 12801
rect 40954 12792 40960 12804
rect 41012 12792 41018 12844
rect 43901 12835 43959 12841
rect 43901 12801 43913 12835
rect 43947 12801 43959 12835
rect 44082 12832 44088 12844
rect 44043 12804 44088 12832
rect 43901 12795 43959 12801
rect 28966 12736 29500 12764
rect 40862 12724 40868 12776
rect 40920 12764 40926 12776
rect 41233 12767 41291 12773
rect 41233 12764 41245 12767
rect 40920 12736 41245 12764
rect 40920 12724 40926 12736
rect 41233 12733 41245 12736
rect 41279 12733 41291 12767
rect 41233 12727 41291 12733
rect 43916 12764 43944 12795
rect 44082 12792 44088 12804
rect 44140 12792 44146 12844
rect 44174 12792 44180 12844
rect 44232 12832 44238 12844
rect 44269 12835 44327 12841
rect 44269 12832 44281 12835
rect 44232 12804 44281 12832
rect 44232 12792 44238 12804
rect 44269 12801 44281 12804
rect 44315 12801 44327 12835
rect 44269 12795 44327 12801
rect 45557 12835 45615 12841
rect 45557 12801 45569 12835
rect 45603 12832 45615 12835
rect 45646 12832 45652 12844
rect 45603 12804 45652 12832
rect 45603 12801 45615 12804
rect 45557 12795 45615 12801
rect 45646 12792 45652 12804
rect 45704 12792 45710 12844
rect 50798 12832 50804 12844
rect 50759 12804 50804 12832
rect 50798 12792 50804 12804
rect 50856 12792 50862 12844
rect 53653 12835 53711 12841
rect 53653 12801 53665 12835
rect 53699 12801 53711 12835
rect 53834 12832 53840 12844
rect 53795 12804 53840 12832
rect 53653 12795 53711 12801
rect 43916 12736 44312 12764
rect 24670 12696 24676 12708
rect 20487 12668 21036 12696
rect 22066 12668 24676 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 17218 12628 17224 12640
rect 16224 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 21008 12637 21036 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 28810 12656 28816 12708
rect 28868 12696 28874 12708
rect 29825 12699 29883 12705
rect 29825 12696 29837 12699
rect 28868 12668 29837 12696
rect 28868 12656 28874 12668
rect 29825 12665 29837 12668
rect 29871 12665 29883 12699
rect 29825 12659 29883 12665
rect 39206 12656 39212 12708
rect 39264 12696 39270 12708
rect 43916 12696 43944 12736
rect 44284 12708 44312 12736
rect 48406 12724 48412 12776
rect 48464 12764 48470 12776
rect 48777 12767 48835 12773
rect 48777 12764 48789 12767
rect 48464 12736 48789 12764
rect 48464 12724 48470 12736
rect 48777 12733 48789 12736
rect 48823 12733 48835 12767
rect 50617 12767 50675 12773
rect 50617 12764 50629 12767
rect 48777 12727 48835 12733
rect 50172 12736 50629 12764
rect 39264 12668 43944 12696
rect 39264 12656 39270 12668
rect 44266 12656 44272 12708
rect 44324 12656 44330 12708
rect 44637 12699 44695 12705
rect 44637 12665 44649 12699
rect 44683 12696 44695 12699
rect 45738 12696 45744 12708
rect 44683 12668 45744 12696
rect 44683 12665 44695 12668
rect 44637 12659 44695 12665
rect 45738 12656 45744 12668
rect 45796 12696 45802 12708
rect 46658 12696 46664 12708
rect 45796 12668 46664 12696
rect 45796 12656 45802 12668
rect 46658 12656 46664 12668
rect 46716 12656 46722 12708
rect 50172 12705 50200 12736
rect 50617 12733 50629 12736
rect 50663 12764 50675 12767
rect 50890 12764 50896 12776
rect 50663 12736 50896 12764
rect 50663 12733 50675 12736
rect 50617 12727 50675 12733
rect 50890 12724 50896 12736
rect 50948 12724 50954 12776
rect 53668 12764 53696 12795
rect 53834 12792 53840 12804
rect 53892 12792 53898 12844
rect 53929 12835 53987 12841
rect 53929 12801 53941 12835
rect 53975 12832 53987 12835
rect 54202 12832 54208 12844
rect 53975 12804 54208 12832
rect 53975 12801 53987 12804
rect 53929 12795 53987 12801
rect 54202 12792 54208 12804
rect 54260 12792 54266 12844
rect 54680 12841 54708 12872
rect 55490 12860 55496 12872
rect 55548 12900 55554 12912
rect 57256 12900 57284 12931
rect 55548 12872 57284 12900
rect 55548 12860 55554 12872
rect 54665 12835 54723 12841
rect 54665 12801 54677 12835
rect 54711 12801 54723 12835
rect 54665 12795 54723 12801
rect 55306 12792 55312 12844
rect 55364 12832 55370 12844
rect 56117 12835 56175 12841
rect 56117 12832 56129 12835
rect 55364 12804 56129 12832
rect 55364 12792 55370 12804
rect 56117 12801 56129 12804
rect 56163 12801 56175 12835
rect 56117 12795 56175 12801
rect 54018 12764 54024 12776
rect 53668 12736 54024 12764
rect 54018 12724 54024 12736
rect 54076 12764 54082 12776
rect 54938 12764 54944 12776
rect 54076 12736 54800 12764
rect 54899 12736 54944 12764
rect 54076 12724 54082 12736
rect 50157 12699 50215 12705
rect 50157 12665 50169 12699
rect 50203 12665 50215 12699
rect 50157 12659 50215 12665
rect 54772 12640 54800 12736
rect 54938 12724 54944 12736
rect 54996 12724 55002 12776
rect 55858 12764 55864 12776
rect 55819 12736 55864 12764
rect 55858 12724 55864 12736
rect 55916 12724 55922 12776
rect 20993 12631 21051 12637
rect 20993 12597 21005 12631
rect 21039 12597 21051 12631
rect 21174 12628 21180 12640
rect 21135 12600 21180 12628
rect 20993 12591 21051 12597
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22554 12628 22560 12640
rect 22152 12600 22560 12628
rect 22152 12588 22158 12600
rect 22554 12588 22560 12600
rect 22612 12628 22618 12640
rect 24213 12631 24271 12637
rect 24213 12628 24225 12631
rect 22612 12600 24225 12628
rect 22612 12588 22618 12600
rect 24213 12597 24225 12600
rect 24259 12597 24271 12631
rect 24213 12591 24271 12597
rect 26142 12588 26148 12640
rect 26200 12628 26206 12640
rect 27430 12628 27436 12640
rect 26200 12600 27436 12628
rect 26200 12588 26206 12600
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 28626 12588 28632 12640
rect 28684 12628 28690 12640
rect 28721 12631 28779 12637
rect 28721 12628 28733 12631
rect 28684 12600 28733 12628
rect 28684 12588 28690 12600
rect 28721 12597 28733 12600
rect 28767 12597 28779 12631
rect 28721 12591 28779 12597
rect 28948 12588 28954 12640
rect 29006 12628 29012 12640
rect 31110 12628 31116 12640
rect 29006 12600 31116 12628
rect 29006 12588 29012 12600
rect 31110 12588 31116 12600
rect 31168 12588 31174 12640
rect 37274 12588 37280 12640
rect 37332 12628 37338 12640
rect 38933 12631 38991 12637
rect 38933 12628 38945 12631
rect 37332 12600 38945 12628
rect 37332 12588 37338 12600
rect 38933 12597 38945 12600
rect 38979 12597 38991 12631
rect 38933 12591 38991 12597
rect 39850 12588 39856 12640
rect 39908 12628 39914 12640
rect 40129 12631 40187 12637
rect 40129 12628 40141 12631
rect 39908 12600 40141 12628
rect 39908 12588 39914 12600
rect 40129 12597 40141 12600
rect 40175 12597 40187 12631
rect 40129 12591 40187 12597
rect 45373 12631 45431 12637
rect 45373 12597 45385 12631
rect 45419 12628 45431 12631
rect 45554 12628 45560 12640
rect 45419 12600 45560 12628
rect 45419 12597 45431 12600
rect 45373 12591 45431 12597
rect 45554 12588 45560 12600
rect 45612 12588 45618 12640
rect 53926 12628 53932 12640
rect 53887 12600 53932 12628
rect 53926 12588 53932 12600
rect 53984 12588 53990 12640
rect 54754 12628 54760 12640
rect 54715 12600 54760 12628
rect 54754 12588 54760 12600
rect 54812 12588 54818 12640
rect 54849 12631 54907 12637
rect 54849 12597 54861 12631
rect 54895 12628 54907 12631
rect 55214 12628 55220 12640
rect 54895 12600 55220 12628
rect 54895 12597 54907 12600
rect 54849 12591 54907 12597
rect 55214 12588 55220 12600
rect 55272 12588 55278 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 2682 12424 2688 12436
rect 2363 12396 2688 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 5902 12424 5908 12436
rect 5863 12396 5908 12424
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 21910 12424 21916 12436
rect 6012 12396 17264 12424
rect 21871 12396 21916 12424
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 6012 12356 6040 12396
rect 4120 12328 6040 12356
rect 4120 12316 4126 12328
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 7524 12328 10057 12356
rect 7524 12316 7530 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2869 12291 2927 12297
rect 2869 12288 2881 12291
rect 2648 12260 2881 12288
rect 2648 12248 2654 12260
rect 2869 12257 2881 12260
rect 2915 12288 2927 12291
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 2915 12260 4445 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 4433 12257 4445 12260
rect 4479 12257 4491 12291
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 4433 12251 4491 12257
rect 6886 12260 9321 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1452 12192 1593 12220
rect 1452 12180 1458 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12220 4307 12223
rect 4614 12220 4620 12232
rect 4295 12192 4620 12220
rect 4295 12189 4307 12192
rect 4249 12183 4307 12189
rect 4614 12180 4620 12192
rect 4672 12220 4678 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 4672 12192 6193 12220
rect 4672 12180 4678 12192
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 2777 12155 2835 12161
rect 2777 12152 2789 12155
rect 1412 12124 2789 12152
rect 1412 12093 1440 12124
rect 2777 12121 2789 12124
rect 2823 12121 2835 12155
rect 2777 12115 2835 12121
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 5537 12155 5595 12161
rect 5537 12152 5549 12155
rect 5500 12124 5549 12152
rect 5500 12112 5506 12124
rect 5537 12121 5549 12124
rect 5583 12152 5595 12155
rect 6886 12152 6914 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 10060 12288 10088 12319
rect 10226 12316 10232 12368
rect 10284 12356 10290 12368
rect 10778 12356 10784 12368
rect 10284 12328 10784 12356
rect 10284 12316 10290 12328
rect 10778 12316 10784 12328
rect 10836 12356 10842 12368
rect 11057 12359 11115 12365
rect 11057 12356 11069 12359
rect 10836 12328 11069 12356
rect 10836 12316 10842 12328
rect 11057 12325 11069 12328
rect 11103 12325 11115 12359
rect 17236 12356 17264 12396
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 32214 12424 32220 12436
rect 22066 12396 32220 12424
rect 22066 12356 22094 12396
rect 32214 12384 32220 12396
rect 32272 12384 32278 12436
rect 32490 12384 32496 12436
rect 32548 12424 32554 12436
rect 32585 12427 32643 12433
rect 32585 12424 32597 12427
rect 32548 12396 32597 12424
rect 32548 12384 32554 12396
rect 32585 12393 32597 12396
rect 32631 12393 32643 12427
rect 34514 12424 34520 12436
rect 32585 12387 32643 12393
rect 33796 12396 34520 12424
rect 22738 12356 22744 12368
rect 17236 12328 22094 12356
rect 22699 12328 22744 12356
rect 11057 12319 11115 12325
rect 22738 12316 22744 12328
rect 22796 12316 22802 12368
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 26605 12359 26663 12365
rect 26605 12356 26617 12359
rect 24176 12328 26617 12356
rect 24176 12316 24182 12328
rect 26605 12325 26617 12328
rect 26651 12325 26663 12359
rect 32232 12356 32260 12384
rect 33321 12359 33379 12365
rect 33321 12356 33333 12359
rect 32232 12328 33333 12356
rect 26605 12319 26663 12325
rect 33321 12325 33333 12328
rect 33367 12325 33379 12359
rect 33321 12319 33379 12325
rect 11606 12288 11612 12300
rect 9456 12260 9501 12288
rect 10060 12260 11612 12288
rect 9456 12248 9462 12260
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 19426 12288 19432 12300
rect 17276 12260 19432 12288
rect 17276 12248 17282 12260
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 21450 12248 21456 12300
rect 21508 12288 21514 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21508 12260 22017 12288
rect 21508 12248 21514 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 27709 12291 27767 12297
rect 27709 12288 27721 12291
rect 22152 12260 27721 12288
rect 22152 12248 22158 12260
rect 27709 12257 27721 12260
rect 27755 12288 27767 12291
rect 28077 12291 28135 12297
rect 28077 12288 28089 12291
rect 27755 12260 28089 12288
rect 27755 12257 27767 12260
rect 27709 12251 27767 12257
rect 28077 12257 28089 12260
rect 28123 12257 28135 12291
rect 28077 12251 28135 12257
rect 7098 12220 7104 12232
rect 7059 12192 7104 12220
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 7248 12192 7297 12220
rect 7248 12180 7254 12192
rect 7285 12189 7297 12192
rect 7331 12220 7343 12223
rect 7742 12220 7748 12232
rect 7331 12192 7748 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 9030 12220 9036 12232
rect 8312 12192 9036 12220
rect 5583 12124 6914 12152
rect 7116 12152 7144 12180
rect 7374 12152 7380 12164
rect 7116 12124 7380 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 7374 12112 7380 12124
rect 7432 12152 7438 12164
rect 8205 12155 8263 12161
rect 8205 12152 8217 12155
rect 7432 12124 8217 12152
rect 7432 12112 7438 12124
rect 8205 12121 8217 12124
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 1397 12087 1455 12093
rect 1397 12053 1409 12087
rect 1443 12053 1455 12087
rect 2682 12084 2688 12096
rect 2643 12056 2688 12084
rect 1397 12047 1455 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 5914 12087 5972 12093
rect 5914 12053 5926 12087
rect 5960 12084 5972 12087
rect 6730 12084 6736 12096
rect 5960 12056 6736 12084
rect 5960 12053 5972 12056
rect 5914 12047 5972 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 8312 12084 8340 12192
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 8389 12155 8447 12161
rect 8389 12121 8401 12155
rect 8435 12152 8447 12155
rect 9140 12152 9168 12183
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9490 12220 9496 12232
rect 9272 12192 9496 12220
rect 9272 12180 9278 12192
rect 9490 12180 9496 12192
rect 9548 12220 9554 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9548 12192 9873 12220
rect 9548 12180 9554 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 10502 12220 10508 12232
rect 9861 12183 9919 12189
rect 10060 12192 10508 12220
rect 10060 12152 10088 12192
rect 10502 12180 10508 12192
rect 10560 12220 10566 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 10560 12192 10701 12220
rect 10560 12180 10566 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10870 12220 10876 12232
rect 10831 12192 10876 12220
rect 10689 12183 10747 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 14332 12192 14473 12220
rect 14332 12180 14338 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 16724 12192 17877 12220
rect 16724 12180 16730 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 18138 12220 18144 12232
rect 18099 12192 18144 12220
rect 17865 12183 17923 12189
rect 18138 12180 18144 12192
rect 18196 12220 18202 12232
rect 18414 12220 18420 12232
rect 18196 12192 18420 12220
rect 18196 12180 18202 12192
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21324 12192 21925 12220
rect 21324 12180 21330 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 22922 12220 22928 12232
rect 22883 12192 22928 12220
rect 21913 12183 21971 12189
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 23014 12180 23020 12232
rect 23072 12220 23078 12232
rect 23072 12192 23117 12220
rect 23072 12180 23078 12192
rect 25314 12180 25320 12232
rect 25372 12220 25378 12232
rect 25961 12223 26019 12229
rect 25961 12220 25973 12223
rect 25372 12192 25973 12220
rect 25372 12180 25378 12192
rect 25961 12189 25973 12192
rect 26007 12189 26019 12223
rect 25961 12183 26019 12189
rect 26054 12223 26112 12229
rect 26054 12189 26066 12223
rect 26100 12220 26112 12223
rect 26142 12220 26148 12232
rect 26100 12192 26148 12220
rect 26100 12189 26112 12192
rect 26054 12183 26112 12189
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 26237 12223 26295 12229
rect 26237 12189 26249 12223
rect 26283 12220 26295 12223
rect 26283 12189 26296 12220
rect 26237 12183 26296 12189
rect 8435 12124 9076 12152
rect 9140 12124 10088 12152
rect 14728 12155 14786 12161
rect 8435 12121 8447 12124
rect 8389 12115 8447 12121
rect 7239 12056 8340 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8904 12056 8953 12084
rect 8904 12044 8910 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 9048 12084 9076 12124
rect 14728 12121 14740 12155
rect 14774 12152 14786 12155
rect 15102 12152 15108 12164
rect 14774 12124 15108 12152
rect 14774 12121 14786 12124
rect 14728 12115 14786 12121
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 22646 12152 22652 12164
rect 15988 12124 22652 12152
rect 15988 12112 15994 12124
rect 22646 12112 22652 12124
rect 22704 12112 22710 12164
rect 22741 12155 22799 12161
rect 22741 12121 22753 12155
rect 22787 12152 22799 12155
rect 23566 12152 23572 12164
rect 22787 12124 23572 12152
rect 22787 12121 22799 12124
rect 22741 12115 22799 12121
rect 23566 12112 23572 12124
rect 23624 12112 23630 12164
rect 9398 12084 9404 12096
rect 9048 12056 9404 12084
rect 8941 12047 8999 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10410 12084 10416 12096
rect 9732 12056 10416 12084
rect 9732 12044 9738 12056
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 15286 12084 15292 12096
rect 13596 12056 15292 12084
rect 13596 12044 13602 12056
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 15841 12087 15899 12093
rect 15841 12084 15853 12087
rect 15344 12056 15853 12084
rect 15344 12044 15350 12056
rect 15841 12053 15853 12056
rect 15887 12053 15899 12087
rect 15841 12047 15899 12053
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 22094 12084 22100 12096
rect 16448 12056 22100 12084
rect 16448 12044 16454 12056
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22281 12087 22339 12093
rect 22281 12053 22293 12087
rect 22327 12084 22339 12087
rect 23014 12084 23020 12096
rect 22327 12056 23020 12084
rect 22327 12053 22339 12056
rect 22281 12047 22339 12053
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 25590 12044 25596 12096
rect 25648 12084 25654 12096
rect 26268 12084 26296 12183
rect 26418 12180 26424 12232
rect 26476 12229 26482 12232
rect 26476 12220 26484 12229
rect 26476 12192 26521 12220
rect 26476 12183 26484 12192
rect 26476 12180 26482 12183
rect 26329 12155 26387 12161
rect 26329 12121 26341 12155
rect 26375 12152 26387 12155
rect 27246 12152 27252 12164
rect 26375 12124 27252 12152
rect 26375 12121 26387 12124
rect 26329 12115 26387 12121
rect 27246 12112 27252 12124
rect 27304 12112 27310 12164
rect 26510 12084 26516 12096
rect 25648 12056 26516 12084
rect 25648 12044 25654 12056
rect 26510 12044 26516 12056
rect 26568 12044 26574 12096
rect 28092 12084 28120 12251
rect 30190 12248 30196 12300
rect 30248 12288 30254 12300
rect 33796 12288 33824 12396
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 36078 12384 36084 12436
rect 36136 12424 36142 12436
rect 39209 12427 39267 12433
rect 39209 12424 39221 12427
rect 36136 12396 39221 12424
rect 36136 12384 36142 12396
rect 39209 12393 39221 12396
rect 39255 12424 39267 12427
rect 40310 12424 40316 12436
rect 39255 12396 40316 12424
rect 39255 12393 39267 12396
rect 39209 12387 39267 12393
rect 40310 12384 40316 12396
rect 40368 12384 40374 12436
rect 44266 12384 44272 12436
rect 44324 12424 44330 12436
rect 46661 12427 46719 12433
rect 46661 12424 46673 12427
rect 44324 12396 46673 12424
rect 44324 12384 44330 12396
rect 46661 12393 46673 12396
rect 46707 12393 46719 12427
rect 46661 12387 46719 12393
rect 48961 12427 49019 12433
rect 48961 12393 48973 12427
rect 49007 12424 49019 12427
rect 49142 12424 49148 12436
rect 49007 12396 49148 12424
rect 49007 12393 49019 12396
rect 48961 12387 49019 12393
rect 49142 12384 49148 12396
rect 49200 12384 49206 12436
rect 50433 12427 50491 12433
rect 50433 12424 50445 12427
rect 50080 12396 50445 12424
rect 40037 12359 40095 12365
rect 40037 12356 40049 12359
rect 30248 12260 33824 12288
rect 33888 12328 40049 12356
rect 30248 12248 30254 12260
rect 28166 12180 28172 12232
rect 28224 12220 28230 12232
rect 28353 12223 28411 12229
rect 28353 12220 28365 12223
rect 28224 12192 28365 12220
rect 28224 12180 28230 12192
rect 28353 12189 28365 12192
rect 28399 12189 28411 12223
rect 28353 12183 28411 12189
rect 31573 12223 31631 12229
rect 31573 12189 31585 12223
rect 31619 12220 31631 12223
rect 32122 12220 32128 12232
rect 31619 12192 32128 12220
rect 31619 12189 31631 12192
rect 31573 12183 31631 12189
rect 32122 12180 32128 12192
rect 32180 12180 32186 12232
rect 32306 12220 32312 12232
rect 32267 12192 32312 12220
rect 32306 12180 32312 12192
rect 32364 12180 32370 12232
rect 32401 12223 32459 12229
rect 32401 12189 32413 12223
rect 32447 12220 32459 12223
rect 33321 12223 33379 12229
rect 33321 12220 33333 12223
rect 32447 12192 33333 12220
rect 32447 12189 32459 12192
rect 32401 12183 32459 12189
rect 33321 12189 33333 12192
rect 33367 12220 33379 12223
rect 33888 12220 33916 12328
rect 35897 12291 35955 12297
rect 35897 12257 35909 12291
rect 35943 12288 35955 12291
rect 35943 12260 36952 12288
rect 35943 12257 35955 12260
rect 35897 12251 35955 12257
rect 33367 12192 33916 12220
rect 33367 12189 33379 12192
rect 33321 12183 33379 12189
rect 33962 12180 33968 12232
rect 34020 12220 34026 12232
rect 35805 12223 35863 12229
rect 35805 12220 35817 12223
rect 34020 12192 35817 12220
rect 34020 12180 34026 12192
rect 35805 12189 35817 12192
rect 35851 12189 35863 12223
rect 35805 12183 35863 12189
rect 36538 12180 36544 12232
rect 36596 12220 36602 12232
rect 36924 12229 36952 12260
rect 37016 12229 37044 12328
rect 40037 12325 40049 12328
rect 40083 12356 40095 12359
rect 43625 12359 43683 12365
rect 40083 12328 41460 12356
rect 40083 12325 40095 12328
rect 40037 12319 40095 12325
rect 38626 12260 39436 12288
rect 36633 12223 36691 12229
rect 36633 12220 36645 12223
rect 36596 12192 36645 12220
rect 36596 12180 36602 12192
rect 36633 12189 36645 12192
rect 36679 12189 36691 12223
rect 36633 12183 36691 12189
rect 36725 12223 36783 12229
rect 36725 12189 36737 12223
rect 36771 12189 36783 12223
rect 36725 12183 36783 12189
rect 36909 12223 36967 12229
rect 36909 12189 36921 12223
rect 36955 12189 36967 12223
rect 36909 12183 36967 12189
rect 37001 12223 37059 12229
rect 37001 12189 37013 12223
rect 37047 12220 37059 12223
rect 37090 12220 37096 12232
rect 37047 12192 37096 12220
rect 37047 12189 37059 12192
rect 37001 12183 37059 12189
rect 31754 12112 31760 12164
rect 31812 12152 31818 12164
rect 34698 12152 34704 12164
rect 31812 12124 31857 12152
rect 33244 12124 34704 12152
rect 31812 12112 31818 12124
rect 33244 12084 33272 12124
rect 34698 12112 34704 12124
rect 34756 12112 34762 12164
rect 36740 12152 36768 12183
rect 37090 12180 37096 12192
rect 37148 12180 37154 12232
rect 37274 12180 37280 12232
rect 37332 12220 37338 12232
rect 37645 12223 37703 12229
rect 37645 12220 37657 12223
rect 37332 12192 37657 12220
rect 37332 12180 37338 12192
rect 37645 12189 37657 12192
rect 37691 12189 37703 12223
rect 37645 12183 37703 12189
rect 37829 12223 37887 12229
rect 37829 12189 37841 12223
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 37921 12223 37979 12229
rect 37921 12189 37933 12223
rect 37967 12220 37979 12223
rect 38626 12220 38654 12260
rect 37967 12192 38654 12220
rect 39117 12223 39175 12229
rect 37967 12189 37979 12192
rect 37921 12183 37979 12189
rect 39117 12189 39129 12223
rect 39163 12189 39175 12223
rect 39117 12183 39175 12189
rect 39301 12223 39359 12229
rect 39301 12189 39313 12223
rect 39347 12189 39359 12223
rect 39408 12220 39436 12260
rect 39850 12220 39856 12232
rect 39908 12229 39914 12232
rect 39408 12192 39856 12220
rect 39301 12183 39359 12189
rect 37844 12152 37872 12183
rect 36372 12124 37872 12152
rect 28092 12056 33272 12084
rect 33686 12044 33692 12096
rect 33744 12084 33750 12096
rect 36372 12084 36400 12124
rect 38470 12112 38476 12164
rect 38528 12152 38534 12164
rect 39132 12152 39160 12183
rect 38528 12124 39160 12152
rect 39316 12152 39344 12183
rect 39850 12180 39856 12192
rect 39908 12220 39917 12229
rect 40678 12220 40684 12232
rect 39908 12192 39953 12220
rect 40639 12192 40684 12220
rect 39908 12183 39917 12192
rect 39908 12180 39914 12183
rect 40678 12180 40684 12192
rect 40736 12180 40742 12232
rect 41432 12220 41460 12328
rect 43625 12325 43637 12359
rect 43671 12356 43683 12359
rect 44174 12356 44180 12368
rect 43671 12328 44180 12356
rect 43671 12325 43683 12328
rect 43625 12319 43683 12325
rect 44174 12316 44180 12328
rect 44232 12316 44238 12368
rect 42426 12248 42432 12300
rect 42484 12288 42490 12300
rect 45281 12291 45339 12297
rect 45281 12288 45293 12291
rect 42484 12260 45293 12288
rect 42484 12248 42490 12260
rect 45281 12257 45293 12260
rect 45327 12257 45339 12291
rect 45281 12251 45339 12257
rect 44910 12220 44916 12232
rect 41432 12192 44916 12220
rect 44910 12180 44916 12192
rect 44968 12180 44974 12232
rect 40862 12152 40868 12164
rect 39316 12124 40868 12152
rect 38528 12112 38534 12124
rect 33744 12056 36400 12084
rect 36449 12087 36507 12093
rect 33744 12044 33750 12056
rect 36449 12053 36461 12087
rect 36495 12084 36507 12087
rect 37366 12084 37372 12096
rect 36495 12056 37372 12084
rect 36495 12053 36507 12056
rect 36449 12047 36507 12053
rect 37366 12044 37372 12056
rect 37424 12044 37430 12096
rect 37458 12044 37464 12096
rect 37516 12084 37522 12096
rect 39132 12084 39160 12124
rect 40862 12112 40868 12124
rect 40920 12112 40926 12164
rect 43254 12112 43260 12164
rect 43312 12152 43318 12164
rect 44266 12152 44272 12164
rect 43312 12124 43852 12152
rect 44227 12124 44272 12152
rect 43312 12112 43318 12124
rect 40773 12087 40831 12093
rect 40773 12084 40785 12087
rect 37516 12056 37561 12084
rect 39132 12056 40785 12084
rect 37516 12044 37522 12056
rect 40773 12053 40785 12056
rect 40819 12053 40831 12087
rect 40773 12047 40831 12053
rect 41138 12044 41144 12096
rect 41196 12084 41202 12096
rect 42426 12084 42432 12096
rect 41196 12056 42432 12084
rect 41196 12044 41202 12056
rect 42426 12044 42432 12056
rect 42484 12044 42490 12096
rect 43714 12084 43720 12096
rect 43675 12056 43720 12084
rect 43714 12044 43720 12056
rect 43772 12044 43778 12096
rect 43824 12084 43852 12124
rect 44266 12112 44272 12124
rect 44324 12112 44330 12164
rect 44358 12084 44364 12096
rect 43824 12056 44364 12084
rect 44358 12044 44364 12056
rect 44416 12044 44422 12096
rect 45296 12084 45324 12251
rect 48590 12248 48596 12300
rect 48648 12288 48654 12300
rect 49053 12291 49111 12297
rect 49053 12288 49065 12291
rect 48648 12260 49065 12288
rect 48648 12248 48654 12260
rect 49053 12257 49065 12260
rect 49099 12257 49111 12291
rect 49053 12251 49111 12257
rect 45554 12229 45560 12232
rect 45548 12183 45560 12229
rect 45612 12220 45618 12232
rect 48777 12223 48835 12229
rect 45612 12192 45648 12220
rect 45554 12180 45560 12183
rect 45612 12180 45618 12192
rect 48777 12189 48789 12223
rect 48823 12189 48835 12223
rect 48777 12183 48835 12189
rect 48869 12223 48927 12229
rect 48869 12189 48881 12223
rect 48915 12220 48927 12223
rect 49694 12220 49700 12232
rect 48915 12192 49700 12220
rect 48915 12189 48927 12192
rect 48869 12183 48927 12189
rect 48792 12152 48820 12183
rect 49694 12180 49700 12192
rect 49752 12180 49758 12232
rect 50080 12152 50108 12396
rect 50433 12393 50445 12396
rect 50479 12393 50491 12427
rect 50614 12424 50620 12436
rect 50575 12396 50620 12424
rect 50433 12387 50491 12393
rect 50448 12356 50476 12387
rect 50614 12384 50620 12396
rect 50672 12424 50678 12436
rect 55306 12424 55312 12436
rect 50672 12396 51074 12424
rect 55267 12396 55312 12424
rect 50672 12384 50678 12396
rect 50890 12356 50896 12368
rect 50448 12328 50896 12356
rect 50890 12316 50896 12328
rect 50948 12316 50954 12368
rect 51046 12356 51074 12396
rect 55306 12384 55312 12396
rect 55364 12384 55370 12436
rect 53742 12356 53748 12368
rect 51046 12328 53748 12356
rect 53742 12316 53748 12328
rect 53800 12316 53806 12368
rect 53834 12316 53840 12368
rect 53892 12316 53898 12368
rect 51445 12291 51503 12297
rect 51445 12257 51457 12291
rect 51491 12288 51503 12291
rect 53852 12288 53880 12316
rect 53929 12291 53987 12297
rect 53929 12288 53941 12291
rect 51491 12260 53941 12288
rect 51491 12257 51503 12260
rect 51445 12251 51503 12257
rect 53929 12257 53941 12260
rect 53975 12257 53987 12291
rect 53929 12251 53987 12257
rect 51629 12223 51687 12229
rect 51629 12189 51641 12223
rect 51675 12220 51687 12223
rect 53742 12220 53748 12232
rect 51675 12192 53604 12220
rect 53703 12192 53748 12220
rect 51675 12189 51687 12192
rect 51629 12183 51687 12189
rect 48792 12124 50108 12152
rect 50154 12112 50160 12164
rect 50212 12152 50218 12164
rect 50249 12155 50307 12161
rect 50249 12152 50261 12155
rect 50212 12124 50261 12152
rect 50212 12112 50218 12124
rect 50249 12121 50261 12124
rect 50295 12152 50307 12155
rect 51721 12155 51779 12161
rect 51721 12152 51733 12155
rect 50295 12124 51733 12152
rect 50295 12121 50307 12124
rect 50249 12115 50307 12121
rect 51721 12121 51733 12124
rect 51767 12121 51779 12155
rect 53576 12152 53604 12192
rect 53742 12180 53748 12192
rect 53800 12180 53806 12232
rect 53837 12223 53895 12229
rect 53837 12189 53849 12223
rect 53883 12189 53895 12223
rect 54018 12220 54024 12232
rect 53979 12192 54024 12220
rect 53837 12183 53895 12189
rect 53852 12152 53880 12183
rect 54018 12180 54024 12192
rect 54076 12220 54082 12232
rect 54202 12220 54208 12232
rect 54076 12192 54208 12220
rect 54076 12180 54082 12192
rect 54202 12180 54208 12192
rect 54260 12180 54266 12232
rect 54754 12180 54760 12232
rect 54812 12220 54818 12232
rect 55585 12223 55643 12229
rect 55585 12220 55597 12223
rect 54812 12192 55597 12220
rect 54812 12180 54818 12192
rect 55585 12189 55597 12192
rect 55631 12189 55643 12223
rect 55585 12183 55643 12189
rect 54110 12152 54116 12164
rect 53576 12124 54116 12152
rect 51721 12115 51779 12121
rect 54110 12112 54116 12124
rect 54168 12112 54174 12164
rect 55214 12112 55220 12164
rect 55272 12152 55278 12164
rect 55309 12155 55367 12161
rect 55309 12152 55321 12155
rect 55272 12124 55321 12152
rect 55272 12112 55278 12124
rect 55309 12121 55321 12124
rect 55355 12121 55367 12155
rect 55490 12152 55496 12164
rect 55451 12124 55496 12152
rect 55309 12115 55367 12121
rect 55490 12112 55496 12124
rect 55548 12112 55554 12164
rect 45554 12084 45560 12096
rect 45296 12056 45560 12084
rect 45554 12044 45560 12056
rect 45612 12044 45618 12096
rect 49694 12044 49700 12096
rect 49752 12084 49758 12096
rect 50459 12087 50517 12093
rect 50459 12084 50471 12087
rect 49752 12056 50471 12084
rect 49752 12044 49758 12056
rect 50459 12053 50471 12056
rect 50505 12084 50517 12087
rect 50798 12084 50804 12096
rect 50505 12056 50804 12084
rect 50505 12053 50517 12056
rect 50459 12047 50517 12053
rect 50798 12044 50804 12056
rect 50856 12044 50862 12096
rect 50982 12044 50988 12096
rect 51040 12084 51046 12096
rect 51813 12087 51871 12093
rect 51813 12084 51825 12087
rect 51040 12056 51825 12084
rect 51040 12044 51046 12056
rect 51813 12053 51825 12056
rect 51859 12053 51871 12087
rect 51994 12084 52000 12096
rect 51955 12056 52000 12084
rect 51813 12047 51871 12053
rect 51994 12044 52000 12056
rect 52052 12044 52058 12096
rect 53558 12084 53564 12096
rect 53519 12056 53564 12084
rect 53558 12044 53564 12056
rect 53616 12044 53622 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 2740 11852 3985 11880
rect 2740 11840 2746 11852
rect 3973 11849 3985 11852
rect 4019 11880 4031 11883
rect 7098 11880 7104 11892
rect 4019 11852 7104 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 8754 11880 8760 11892
rect 7239 11852 8760 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 13814 11880 13820 11892
rect 8895 11852 13820 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15102 11880 15108 11892
rect 15063 11852 15108 11880
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 20346 11880 20352 11892
rect 15436 11852 20352 11880
rect 15436 11840 15442 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21091 11883 21149 11889
rect 21091 11849 21103 11883
rect 21137 11880 21149 11883
rect 21266 11880 21272 11892
rect 21137 11852 21272 11880
rect 21137 11849 21149 11852
rect 21091 11843 21149 11849
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 25958 11880 25964 11892
rect 25372 11852 25820 11880
rect 25919 11852 25964 11880
rect 25372 11840 25378 11852
rect 3786 11812 3792 11824
rect 2608 11784 3792 11812
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 2608 11753 2636 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 7466 11812 7472 11824
rect 6788 11784 7472 11812
rect 6788 11772 6794 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 11885 11815 11943 11821
rect 7708 11784 8708 11812
rect 7708 11772 7714 11784
rect 2866 11753 2872 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2096 11716 2605 11744
rect 2096 11704 2102 11716
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2860 11744 2872 11753
rect 2827 11716 2872 11744
rect 2593 11707 2651 11713
rect 2860 11707 2872 11716
rect 2866 11704 2872 11707
rect 2924 11704 2930 11756
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6328 11716 7021 11744
rect 6328 11704 6334 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 7248 11716 7389 11744
rect 7248 11704 7254 11716
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7558 11744 7564 11756
rect 7519 11716 7564 11744
rect 7377 11707 7435 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 8680 11753 8708 11784
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 13538 11812 13544 11824
rect 11931 11784 13544 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 22088 11815 22146 11821
rect 13780 11784 22048 11812
rect 13780 11772 13786 11784
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 8754 11744 8760 11756
rect 8711 11716 8760 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7834 11676 7840 11688
rect 6972 11648 7840 11676
rect 6972 11636 6978 11648
rect 7834 11636 7840 11648
rect 7892 11676 7898 11688
rect 8220 11676 8248 11707
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 10134 11744 10140 11756
rect 10095 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10502 11744 10508 11756
rect 10367 11716 10508 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10652 11716 11529 11744
rect 10652 11704 10658 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11610 11747 11668 11753
rect 11610 11713 11622 11747
rect 11656 11713 11668 11747
rect 11790 11744 11796 11756
rect 11751 11716 11796 11744
rect 11610 11707 11668 11713
rect 7892 11648 8248 11676
rect 8573 11679 8631 11685
rect 7892 11636 7898 11648
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 8619 11648 10241 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 11624 11676 11652 11707
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11974 11704 11980 11756
rect 12032 11753 12038 11756
rect 12032 11744 12040 11753
rect 12032 11716 12077 11744
rect 12032 11707 12040 11716
rect 12032 11704 12038 11707
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 12584 11716 13645 11744
rect 12584 11704 12590 11716
rect 13633 11713 13645 11716
rect 13679 11734 13691 11747
rect 13740 11734 15240 11744
rect 13679 11716 15240 11734
rect 13679 11713 13768 11716
rect 13633 11707 13768 11713
rect 13648 11706 13768 11707
rect 12618 11676 12624 11688
rect 11624 11648 12624 11676
rect 10229 11639 10287 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 13814 11676 13820 11688
rect 13775 11648 13820 11676
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 15212 11676 15240 11716
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15565 11747 15623 11753
rect 15344 11716 15389 11744
rect 15344 11704 15350 11716
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15654 11744 15660 11756
rect 15611 11716 15660 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 18138 11744 18144 11756
rect 17635 11716 18144 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11744 18567 11747
rect 18598 11744 18604 11756
rect 18555 11716 18604 11744
rect 18555 11713 18567 11716
rect 18509 11707 18567 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20956 11716 21005 11744
rect 20956 11704 20962 11716
rect 20993 11713 21005 11716
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 21177 11747 21235 11753
rect 21177 11713 21189 11747
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21450 11744 21456 11756
rect 21315 11716 21456 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15212 11648 15393 11676
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 15473 11679 15531 11685
rect 15473 11645 15485 11679
rect 15519 11676 15531 11679
rect 15746 11676 15752 11688
rect 15519 11648 15752 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 17402 11676 17408 11688
rect 17363 11648 17408 11676
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11645 17555 11679
rect 17678 11676 17684 11688
rect 17639 11648 17684 11676
rect 17497 11639 17555 11645
rect 5350 11568 5356 11620
rect 5408 11608 5414 11620
rect 17221 11611 17279 11617
rect 17221 11608 17233 11611
rect 5408 11580 17233 11608
rect 5408 11568 5414 11580
rect 17221 11577 17233 11580
rect 17267 11577 17279 11611
rect 17221 11571 17279 11577
rect 1397 11543 1455 11549
rect 1397 11509 1409 11543
rect 1443 11540 1455 11543
rect 2498 11540 2504 11552
rect 1443 11512 2504 11540
rect 1443 11509 1455 11512
rect 1397 11503 1455 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6512 11512 7389 11540
rect 6512 11500 6518 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 7377 11503 7435 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 10468 11512 12173 11540
rect 10468 11500 10474 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11540 13323 11543
rect 17310 11540 17316 11552
rect 13311 11512 17316 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17512 11540 17540 11639
rect 17678 11636 17684 11648
rect 17736 11636 17742 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18230 11676 18236 11688
rect 18012 11648 18236 11676
rect 18012 11636 18018 11648
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 21192 11676 21220 11707
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 21818 11744 21824 11756
rect 21779 11716 21824 11744
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 22020 11744 22048 11784
rect 22088 11781 22100 11815
rect 22134 11812 22146 11815
rect 22738 11812 22744 11824
rect 22134 11784 22744 11812
rect 22134 11781 22146 11784
rect 22088 11775 22146 11781
rect 22738 11772 22744 11784
rect 22796 11772 22802 11824
rect 25222 11812 25228 11824
rect 22940 11784 25228 11812
rect 22940 11744 22968 11784
rect 25222 11772 25228 11784
rect 25280 11772 25286 11824
rect 25590 11812 25596 11824
rect 25551 11784 25596 11812
rect 25590 11772 25596 11784
rect 25648 11772 25654 11824
rect 25792 11812 25820 11852
rect 25958 11840 25964 11852
rect 26016 11840 26022 11892
rect 26050 11840 26056 11892
rect 26108 11880 26114 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 26108 11852 27353 11880
rect 26108 11840 26114 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 27525 11883 27583 11889
rect 27525 11849 27537 11883
rect 27571 11880 27583 11883
rect 30466 11880 30472 11892
rect 27571 11852 30472 11880
rect 27571 11849 27583 11852
rect 27525 11843 27583 11849
rect 30466 11840 30472 11852
rect 30524 11840 30530 11892
rect 53377 11883 53435 11889
rect 53377 11880 53389 11883
rect 30576 11852 53389 11880
rect 28074 11812 28080 11824
rect 25792 11784 28080 11812
rect 28074 11772 28080 11784
rect 28132 11772 28138 11824
rect 29914 11812 29920 11824
rect 29875 11784 29920 11812
rect 29914 11772 29920 11784
rect 29972 11772 29978 11824
rect 22020 11716 22968 11744
rect 23014 11704 23020 11756
rect 23072 11744 23078 11756
rect 25314 11744 25320 11756
rect 23072 11716 25320 11744
rect 23072 11704 23078 11716
rect 25314 11704 25320 11716
rect 25372 11704 25378 11756
rect 25465 11747 25523 11753
rect 25465 11713 25477 11747
rect 25511 11744 25523 11747
rect 25682 11744 25688 11756
rect 25511 11713 25544 11744
rect 25643 11716 25688 11744
rect 25465 11707 25544 11713
rect 21634 11676 21640 11688
rect 21192 11648 21640 11676
rect 17586 11568 17592 11620
rect 17644 11608 17650 11620
rect 21192 11608 21220 11648
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 25516 11676 25544 11707
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 25774 11704 25780 11756
rect 25832 11753 25838 11756
rect 25832 11744 25840 11753
rect 25832 11716 25877 11744
rect 25832 11707 25840 11716
rect 25832 11704 25838 11707
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26200 11716 26985 11744
rect 26200 11704 26206 11716
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11744 27307 11747
rect 27338 11744 27344 11756
rect 27295 11716 27344 11744
rect 27295 11713 27307 11716
rect 27249 11707 27307 11713
rect 27172 11676 27200 11707
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 27430 11704 27436 11756
rect 27488 11744 27494 11756
rect 30576 11744 30604 11852
rect 53377 11849 53389 11852
rect 53423 11849 53435 11883
rect 53377 11843 53435 11849
rect 30650 11772 30656 11824
rect 30708 11812 30714 11824
rect 33962 11812 33968 11824
rect 30708 11784 33968 11812
rect 30708 11772 30714 11784
rect 33962 11772 33968 11784
rect 34020 11772 34026 11824
rect 34181 11815 34239 11821
rect 34181 11781 34193 11815
rect 34227 11812 34239 11815
rect 35986 11812 35992 11824
rect 34227 11784 35992 11812
rect 34227 11781 34239 11784
rect 34181 11775 34239 11781
rect 35986 11772 35992 11784
rect 36044 11772 36050 11824
rect 37277 11815 37335 11821
rect 37277 11812 37289 11815
rect 36188 11784 37289 11812
rect 32122 11744 32128 11756
rect 27488 11716 30604 11744
rect 32083 11716 32128 11744
rect 27488 11704 27494 11716
rect 32122 11704 32128 11716
rect 32180 11704 32186 11756
rect 34514 11704 34520 11756
rect 34572 11744 34578 11756
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 34572 11716 34805 11744
rect 34572 11704 34578 11716
rect 34793 11713 34805 11716
rect 34839 11713 34851 11747
rect 34793 11707 34851 11713
rect 35060 11747 35118 11753
rect 35060 11713 35072 11747
rect 35106 11744 35118 11747
rect 35342 11744 35348 11756
rect 35106 11716 35348 11744
rect 35106 11713 35118 11716
rect 35060 11707 35118 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 28534 11676 28540 11688
rect 23216 11648 27200 11676
rect 28495 11648 28540 11676
rect 23216 11620 23244 11648
rect 28534 11636 28540 11648
rect 28592 11636 28598 11688
rect 28813 11679 28871 11685
rect 28813 11645 28825 11679
rect 28859 11645 28871 11679
rect 28813 11639 28871 11645
rect 23198 11608 23204 11620
rect 17644 11580 21220 11608
rect 23111 11580 23204 11608
rect 17644 11568 17650 11580
rect 23198 11568 23204 11580
rect 23256 11568 23262 11620
rect 23290 11568 23296 11620
rect 23348 11608 23354 11620
rect 26050 11608 26056 11620
rect 23348 11580 26056 11608
rect 23348 11568 23354 11580
rect 26050 11568 26056 11580
rect 26108 11568 26114 11620
rect 28718 11608 28724 11620
rect 26436 11580 28724 11608
rect 26436 11552 26464 11580
rect 28718 11568 28724 11580
rect 28776 11608 28782 11620
rect 28828 11608 28856 11639
rect 32306 11636 32312 11688
rect 32364 11676 32370 11688
rect 32401 11679 32459 11685
rect 32401 11676 32413 11679
rect 32364 11648 32413 11676
rect 32364 11636 32370 11648
rect 32401 11645 32413 11648
rect 32447 11645 32459 11679
rect 32401 11639 32459 11645
rect 36188 11617 36216 11784
rect 37277 11781 37289 11784
rect 37323 11781 37335 11815
rect 37277 11775 37335 11781
rect 37366 11772 37372 11824
rect 37424 11812 37430 11824
rect 37493 11815 37551 11821
rect 37493 11812 37505 11815
rect 37424 11784 37505 11812
rect 37424 11772 37430 11784
rect 37493 11781 37505 11784
rect 37539 11812 37551 11815
rect 44729 11815 44787 11821
rect 37539 11784 40632 11812
rect 37539 11781 37551 11784
rect 37493 11775 37551 11781
rect 37090 11704 37096 11756
rect 37148 11744 37154 11756
rect 38289 11747 38347 11753
rect 38289 11744 38301 11747
rect 37148 11716 38301 11744
rect 37148 11704 37154 11716
rect 38289 11713 38301 11716
rect 38335 11713 38347 11747
rect 38289 11707 38347 11713
rect 38565 11747 38623 11753
rect 38565 11713 38577 11747
rect 38611 11713 38623 11747
rect 39206 11744 39212 11756
rect 39167 11716 39212 11744
rect 38565 11707 38623 11713
rect 38378 11636 38384 11688
rect 38436 11636 38442 11688
rect 38580 11676 38608 11707
rect 39206 11704 39212 11716
rect 39264 11704 39270 11756
rect 39301 11747 39359 11753
rect 39301 11713 39313 11747
rect 39347 11744 39359 11747
rect 39850 11744 39856 11756
rect 39347 11716 39856 11744
rect 39347 11713 39359 11716
rect 39301 11707 39359 11713
rect 39850 11704 39856 11716
rect 39908 11704 39914 11756
rect 40218 11744 40224 11756
rect 40179 11716 40224 11744
rect 40218 11704 40224 11716
rect 40276 11704 40282 11756
rect 40310 11704 40316 11756
rect 40368 11744 40374 11756
rect 40604 11753 40632 11784
rect 44729 11781 44741 11815
rect 44775 11812 44787 11815
rect 44818 11812 44824 11824
rect 44775 11784 44824 11812
rect 44775 11781 44787 11784
rect 44729 11775 44787 11781
rect 44818 11772 44824 11784
rect 44876 11772 44882 11824
rect 44945 11815 45003 11821
rect 44945 11781 44957 11815
rect 44991 11812 45003 11815
rect 45738 11812 45744 11824
rect 44991 11784 45744 11812
rect 44991 11781 45003 11784
rect 44945 11775 45003 11781
rect 45738 11772 45744 11784
rect 45796 11772 45802 11824
rect 48498 11812 48504 11824
rect 48459 11784 48504 11812
rect 48498 11772 48504 11784
rect 48556 11772 48562 11824
rect 51445 11815 51503 11821
rect 51445 11781 51457 11815
rect 51491 11781 51503 11815
rect 51445 11775 51503 11781
rect 41248 11753 41392 11766
rect 40589 11747 40647 11753
rect 40368 11716 40413 11744
rect 40368 11704 40374 11716
rect 40589 11713 40601 11747
rect 40635 11713 40647 11747
rect 41248 11747 41429 11753
rect 41248 11744 41383 11747
rect 40589 11707 40647 11713
rect 41064 11738 41383 11744
rect 41064 11716 41276 11738
rect 41364 11716 41383 11738
rect 39224 11676 39252 11704
rect 41064 11688 41092 11716
rect 41371 11713 41383 11716
rect 41417 11713 41429 11747
rect 41371 11707 41429 11713
rect 41487 11704 41493 11756
rect 41545 11753 41551 11756
rect 41545 11747 41564 11753
rect 41552 11713 41564 11747
rect 41545 11707 41564 11713
rect 41601 11747 41659 11753
rect 41601 11713 41613 11747
rect 41647 11713 41659 11747
rect 41601 11707 41659 11713
rect 41797 11747 41855 11753
rect 41966 11747 41972 11756
rect 41797 11713 41809 11747
rect 41843 11719 41972 11747
rect 41843 11713 41855 11719
rect 41797 11707 41855 11713
rect 41545 11704 41551 11707
rect 38580 11648 39252 11676
rect 40497 11679 40555 11685
rect 40497 11645 40509 11679
rect 40543 11676 40555 11679
rect 41046 11676 41052 11688
rect 40543 11648 41052 11676
rect 40543 11645 40555 11648
rect 40497 11639 40555 11645
rect 41046 11636 41052 11648
rect 41104 11636 41110 11688
rect 41138 11636 41144 11688
rect 41196 11676 41202 11688
rect 41196 11648 41241 11676
rect 41196 11636 41202 11648
rect 36173 11611 36231 11617
rect 28776 11580 28856 11608
rect 32232 11580 34192 11608
rect 28776 11568 28782 11580
rect 32232 11552 32260 11580
rect 23106 11540 23112 11552
rect 17512 11512 23112 11540
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 25774 11500 25780 11552
rect 25832 11540 25838 11552
rect 26418 11540 26424 11552
rect 25832 11512 26424 11540
rect 25832 11500 25838 11512
rect 26418 11500 26424 11512
rect 26476 11500 26482 11552
rect 30193 11543 30251 11549
rect 30193 11509 30205 11543
rect 30239 11540 30251 11543
rect 30282 11540 30288 11552
rect 30239 11512 30288 11540
rect 30239 11509 30251 11512
rect 30193 11503 30251 11509
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 32214 11540 32220 11552
rect 32175 11512 32220 11540
rect 32214 11500 32220 11512
rect 32272 11500 32278 11552
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 32950 11540 32956 11552
rect 32355 11512 32956 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 32950 11500 32956 11512
rect 33008 11500 33014 11552
rect 33318 11500 33324 11552
rect 33376 11540 33382 11552
rect 33870 11540 33876 11552
rect 33376 11512 33876 11540
rect 33376 11500 33382 11512
rect 33870 11500 33876 11512
rect 33928 11500 33934 11552
rect 34164 11549 34192 11580
rect 36173 11577 36185 11611
rect 36219 11608 36231 11611
rect 36354 11608 36360 11620
rect 36219 11580 36360 11608
rect 36219 11577 36231 11580
rect 36173 11571 36231 11577
rect 36354 11568 36360 11580
rect 36412 11568 36418 11620
rect 38396 11608 38424 11636
rect 39485 11611 39543 11617
rect 39485 11608 39497 11611
rect 38396 11580 39497 11608
rect 39485 11577 39497 11580
rect 39531 11577 39543 11611
rect 39485 11571 39543 11577
rect 40681 11611 40739 11617
rect 40681 11577 40693 11611
rect 40727 11608 40739 11611
rect 41616 11608 41644 11707
rect 41966 11704 41972 11719
rect 42024 11704 42030 11756
rect 42518 11704 42524 11756
rect 42576 11744 42582 11756
rect 42685 11747 42743 11753
rect 42685 11744 42697 11747
rect 42576 11716 42697 11744
rect 42576 11704 42582 11716
rect 42685 11713 42697 11716
rect 42731 11713 42743 11747
rect 42685 11707 42743 11713
rect 48133 11747 48191 11753
rect 48133 11713 48145 11747
rect 48179 11744 48191 11747
rect 49694 11744 49700 11756
rect 48179 11716 49700 11744
rect 48179 11713 48191 11716
rect 48133 11707 48191 11713
rect 49694 11704 49700 11716
rect 49752 11704 49758 11756
rect 51460 11744 51488 11775
rect 51534 11772 51540 11824
rect 51592 11812 51598 11824
rect 51645 11815 51703 11821
rect 51645 11812 51657 11815
rect 51592 11784 51657 11812
rect 51592 11772 51598 11784
rect 51645 11781 51657 11784
rect 51691 11781 51703 11815
rect 53392 11812 53420 11843
rect 53558 11840 53564 11892
rect 53616 11880 53622 11892
rect 53945 11883 54003 11889
rect 53945 11880 53957 11883
rect 53616 11852 53957 11880
rect 53616 11840 53622 11852
rect 53945 11849 53957 11852
rect 53991 11849 54003 11883
rect 53945 11843 54003 11849
rect 54113 11883 54171 11889
rect 54113 11849 54125 11883
rect 54159 11849 54171 11883
rect 54113 11843 54171 11849
rect 55217 11883 55275 11889
rect 55217 11849 55229 11883
rect 55263 11849 55275 11883
rect 55217 11843 55275 11849
rect 53650 11812 53656 11824
rect 53392 11784 53656 11812
rect 51645 11775 51703 11781
rect 53650 11772 53656 11784
rect 53708 11812 53714 11824
rect 53745 11815 53803 11821
rect 53745 11812 53757 11815
rect 53708 11784 53757 11812
rect 53708 11772 53714 11784
rect 53745 11781 53757 11784
rect 53791 11781 53803 11815
rect 53745 11775 53803 11781
rect 54018 11744 54024 11756
rect 51460 11716 54024 11744
rect 54018 11704 54024 11716
rect 54076 11704 54082 11756
rect 54128 11744 54156 11843
rect 55232 11812 55260 11843
rect 56106 11815 56164 11821
rect 56106 11812 56118 11815
rect 55232 11784 56118 11812
rect 56106 11781 56118 11784
rect 56152 11781 56164 11815
rect 56106 11775 56164 11781
rect 55401 11747 55459 11753
rect 55401 11744 55413 11747
rect 54128 11716 55413 11744
rect 55401 11713 55413 11716
rect 55447 11713 55459 11747
rect 55858 11744 55864 11756
rect 55819 11716 55864 11744
rect 55401 11707 55459 11713
rect 55858 11704 55864 11716
rect 55916 11704 55922 11756
rect 42426 11676 42432 11688
rect 42387 11648 42432 11676
rect 42426 11636 42432 11648
rect 42484 11636 42490 11688
rect 40727 11580 41644 11608
rect 43809 11611 43867 11617
rect 40727 11577 40739 11580
rect 40681 11571 40739 11577
rect 43809 11577 43821 11611
rect 43855 11608 43867 11611
rect 44082 11608 44088 11620
rect 43855 11580 44088 11608
rect 43855 11577 43867 11580
rect 43809 11571 43867 11577
rect 44082 11568 44088 11580
rect 44140 11568 44146 11620
rect 45097 11611 45155 11617
rect 45097 11577 45109 11611
rect 45143 11608 45155 11611
rect 45646 11608 45652 11620
rect 45143 11580 45652 11608
rect 45143 11577 45155 11580
rect 45097 11571 45155 11577
rect 45646 11568 45652 11580
rect 45704 11568 45710 11620
rect 51994 11608 52000 11620
rect 51644 11580 52000 11608
rect 34149 11543 34207 11549
rect 34149 11509 34161 11543
rect 34195 11509 34207 11543
rect 34149 11503 34207 11509
rect 34333 11543 34391 11549
rect 34333 11509 34345 11543
rect 34379 11540 34391 11543
rect 35526 11540 35532 11552
rect 34379 11512 35532 11540
rect 34379 11509 34391 11512
rect 34333 11503 34391 11509
rect 35526 11500 35532 11512
rect 35584 11500 35590 11552
rect 36078 11500 36084 11552
rect 36136 11540 36142 11552
rect 37461 11543 37519 11549
rect 37461 11540 37473 11543
rect 36136 11512 37473 11540
rect 36136 11500 36142 11512
rect 37461 11509 37473 11512
rect 37507 11509 37519 11543
rect 37461 11503 37519 11509
rect 37550 11500 37556 11552
rect 37608 11540 37614 11552
rect 37645 11543 37703 11549
rect 37645 11540 37657 11543
rect 37608 11512 37657 11540
rect 37608 11500 37614 11512
rect 37645 11509 37657 11512
rect 37691 11509 37703 11543
rect 37645 11503 37703 11509
rect 37734 11500 37740 11552
rect 37792 11540 37798 11552
rect 38381 11543 38439 11549
rect 38381 11540 38393 11543
rect 37792 11512 38393 11540
rect 37792 11500 37798 11512
rect 38381 11509 38393 11512
rect 38427 11509 38439 11543
rect 44910 11540 44916 11552
rect 44871 11512 44916 11540
rect 38381 11503 38439 11509
rect 44910 11500 44916 11512
rect 44968 11500 44974 11552
rect 48222 11500 48228 11552
rect 48280 11540 48286 11552
rect 48501 11543 48559 11549
rect 48501 11540 48513 11543
rect 48280 11512 48513 11540
rect 48280 11500 48286 11512
rect 48501 11509 48513 11512
rect 48547 11509 48559 11543
rect 48501 11503 48559 11509
rect 48590 11500 48596 11552
rect 48648 11540 48654 11552
rect 51644 11549 51672 11580
rect 51994 11568 52000 11580
rect 52052 11568 52058 11620
rect 54036 11608 54064 11704
rect 54036 11580 55352 11608
rect 48685 11543 48743 11549
rect 48685 11540 48697 11543
rect 48648 11512 48697 11540
rect 48648 11500 48654 11512
rect 48685 11509 48697 11512
rect 48731 11509 48743 11543
rect 48685 11503 48743 11509
rect 51629 11543 51687 11549
rect 51629 11509 51641 11543
rect 51675 11509 51687 11543
rect 51810 11540 51816 11552
rect 51771 11512 51816 11540
rect 51629 11503 51687 11509
rect 51810 11500 51816 11512
rect 51868 11500 51874 11552
rect 53926 11540 53932 11552
rect 53887 11512 53932 11540
rect 53926 11500 53932 11512
rect 53984 11500 53990 11552
rect 55324 11540 55352 11580
rect 57241 11543 57299 11549
rect 57241 11540 57253 11543
rect 55324 11512 57253 11540
rect 57241 11509 57253 11512
rect 57287 11509 57299 11543
rect 57241 11503 57299 11509
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 10594 11336 10600 11348
rect 10555 11308 10600 11336
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 11848 11308 12357 11336
rect 11848 11296 11854 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 15528 11308 16221 11336
rect 15528 11296 15534 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 17460 11308 18061 11336
rect 17460 11296 17466 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 19260 11308 20300 11336
rect 1578 11268 1584 11280
rect 1539 11240 1584 11268
rect 1578 11228 1584 11240
rect 1636 11228 1642 11280
rect 6822 11228 6828 11280
rect 6880 11268 6886 11280
rect 7190 11268 7196 11280
rect 6880 11240 7196 11268
rect 6880 11228 6886 11240
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 9766 11228 9772 11280
rect 9824 11268 9830 11280
rect 11054 11268 11060 11280
rect 9824 11240 11060 11268
rect 9824 11228 9830 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11606 11268 11612 11280
rect 11567 11240 11612 11268
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 16393 11271 16451 11277
rect 16393 11268 16405 11271
rect 15488 11240 16405 11268
rect 4062 11200 4068 11212
rect 1412 11172 4068 11200
rect 1412 11141 1440 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 7006 11200 7012 11212
rect 6503 11172 7012 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 7006 11160 7012 11172
rect 7064 11200 7070 11212
rect 7558 11200 7564 11212
rect 7064 11172 7564 11200
rect 7064 11160 7070 11172
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 15194 11200 15200 11212
rect 15155 11172 15200 11200
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 15488 11209 15516 11240
rect 16393 11237 16405 11240
rect 16439 11237 16451 11271
rect 16393 11231 16451 11237
rect 17310 11228 17316 11280
rect 17368 11268 17374 11280
rect 19260 11268 19288 11308
rect 17368 11240 19288 11268
rect 17368 11228 17374 11240
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 18046 11160 18052 11212
rect 18104 11200 18110 11212
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 18104 11172 18245 11200
rect 18104 11160 18110 11172
rect 18233 11169 18245 11172
rect 18279 11169 18291 11203
rect 18233 11163 18291 11169
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18509 11203 18567 11209
rect 18380 11172 18425 11200
rect 18380 11160 18386 11172
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 18598 11200 18604 11212
rect 18555 11172 18604 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 20272 11200 20300 11308
rect 20898 11296 20904 11348
rect 20956 11336 20962 11348
rect 20956 11308 22324 11336
rect 20956 11296 20962 11308
rect 22296 11280 22324 11308
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 22554 11336 22560 11348
rect 22428 11308 22473 11336
rect 22515 11308 22560 11336
rect 22428 11296 22434 11308
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 23106 11296 23112 11348
rect 23164 11336 23170 11348
rect 23845 11339 23903 11345
rect 23845 11336 23857 11339
rect 23164 11308 23857 11336
rect 23164 11296 23170 11308
rect 23845 11305 23857 11308
rect 23891 11305 23903 11339
rect 23845 11299 23903 11305
rect 25222 11296 25228 11348
rect 25280 11336 25286 11348
rect 27709 11339 27767 11345
rect 27709 11336 27721 11339
rect 25280 11308 27721 11336
rect 25280 11296 25286 11308
rect 27709 11305 27721 11308
rect 27755 11336 27767 11339
rect 30650 11336 30656 11348
rect 27755 11308 30656 11336
rect 27755 11305 27767 11308
rect 27709 11299 27767 11305
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 32306 11296 32312 11348
rect 32364 11336 32370 11348
rect 32493 11339 32551 11345
rect 32493 11336 32505 11339
rect 32364 11308 32505 11336
rect 32364 11296 32370 11308
rect 32493 11305 32505 11308
rect 32539 11305 32551 11339
rect 32493 11299 32551 11305
rect 33321 11339 33379 11345
rect 33321 11305 33333 11339
rect 33367 11336 33379 11339
rect 33594 11336 33600 11348
rect 33367 11308 33600 11336
rect 33367 11305 33379 11308
rect 33321 11299 33379 11305
rect 33594 11296 33600 11308
rect 33652 11296 33658 11348
rect 35161 11339 35219 11345
rect 35161 11305 35173 11339
rect 35207 11336 35219 11339
rect 35342 11336 35348 11348
rect 35207 11308 35348 11336
rect 35207 11305 35219 11308
rect 35161 11299 35219 11305
rect 35342 11296 35348 11308
rect 35400 11296 35406 11348
rect 35526 11336 35532 11348
rect 35487 11308 35532 11336
rect 35526 11296 35532 11308
rect 35584 11296 35590 11348
rect 35710 11296 35716 11348
rect 35768 11336 35774 11348
rect 38746 11336 38752 11348
rect 35768 11308 38752 11336
rect 35768 11296 35774 11308
rect 38746 11296 38752 11308
rect 38804 11296 38810 11348
rect 40218 11296 40224 11348
rect 40276 11336 40282 11348
rect 47670 11336 47676 11348
rect 40276 11308 47676 11336
rect 40276 11296 40282 11308
rect 47670 11296 47676 11308
rect 47728 11296 47734 11348
rect 48590 11336 48596 11348
rect 47780 11308 48596 11336
rect 20346 11228 20352 11280
rect 20404 11268 20410 11280
rect 22186 11268 22192 11280
rect 20404 11240 22192 11268
rect 20404 11228 20410 11240
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 23198 11268 23204 11280
rect 22336 11240 23204 11268
rect 22336 11228 22342 11240
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 25409 11271 25467 11277
rect 25409 11237 25421 11271
rect 25455 11237 25467 11271
rect 25409 11231 25467 11237
rect 25424 11200 25452 11231
rect 25498 11228 25504 11280
rect 25556 11268 25562 11280
rect 26142 11268 26148 11280
rect 25556 11240 26148 11268
rect 25556 11228 25562 11240
rect 26142 11228 26148 11240
rect 26200 11228 26206 11280
rect 33413 11271 33471 11277
rect 33413 11237 33425 11271
rect 33459 11237 33471 11271
rect 43254 11268 43260 11280
rect 33413 11231 33471 11237
rect 33520 11240 43260 11268
rect 20272 11172 24624 11200
rect 25424 11172 26464 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 1397 11095 1455 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6178 11132 6184 11144
rect 6135 11104 6184 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6362 11132 6368 11144
rect 6323 11104 6368 11132
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6914 11132 6920 11144
rect 6687 11104 6920 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7190 11132 7196 11144
rect 7147 11104 7196 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7374 11132 7380 11144
rect 7335 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11103 11104 11652 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 9950 11064 9956 11076
rect 2884 11036 9956 11064
rect 2225 10999 2283 11005
rect 2225 10965 2237 10999
rect 2271 10996 2283 10999
rect 2314 10996 2320 11008
rect 2271 10968 2320 10996
rect 2271 10965 2283 10968
rect 2225 10959 2283 10965
rect 2314 10956 2320 10968
rect 2372 10956 2378 11008
rect 2884 11005 2912 11036
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 11624 11073 11652 11104
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12342 11132 12348 11144
rect 12207 11104 12348 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11132 15439 11135
rect 15746 11132 15752 11144
rect 15427 11104 15752 11132
rect 15427 11101 15439 11104
rect 15381 11095 15439 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 18414 11132 18420 11144
rect 15856 11104 16344 11132
rect 18375 11104 18420 11132
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 10100 11036 10977 11064
rect 10100 11024 10106 11036
rect 10965 11033 10977 11036
rect 11011 11033 11023 11067
rect 10965 11027 11023 11033
rect 11609 11067 11667 11073
rect 11609 11033 11621 11067
rect 11655 11064 11667 11067
rect 12084 11064 12112 11092
rect 13722 11064 13728 11076
rect 11655 11036 12112 11064
rect 12176 11036 13728 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10965 2927 10999
rect 2869 10959 2927 10965
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11146 10996 11152 11008
rect 10836 10968 11152 10996
rect 10836 10956 10842 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 12069 10999 12127 11005
rect 12069 10965 12081 10999
rect 12115 10996 12127 10999
rect 12176 10996 12204 11036
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 14366 11024 14372 11076
rect 14424 11064 14430 11076
rect 15856 11064 15884 11104
rect 16022 11064 16028 11076
rect 14424 11036 15884 11064
rect 15983 11036 16028 11064
rect 14424 11024 14430 11036
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 16225 11067 16283 11073
rect 16225 11064 16237 11067
rect 16172 11036 16237 11064
rect 16172 11024 16178 11036
rect 16225 11033 16237 11036
rect 16271 11033 16283 11067
rect 16316 11064 16344 11104
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 21376 11104 22784 11132
rect 19518 11073 19524 11076
rect 16316 11036 19334 11064
rect 16225 11027 16283 11033
rect 15010 10996 15016 11008
rect 12115 10968 12204 10996
rect 14971 10968 15016 10996
rect 12115 10965 12127 10968
rect 12069 10959 12127 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 19306 10996 19334 11036
rect 19512 11027 19524 11073
rect 19576 11064 19582 11076
rect 21376 11064 21404 11104
rect 19576 11036 19612 11064
rect 19720 11036 21404 11064
rect 19518 11024 19524 11027
rect 19576 11024 19582 11036
rect 19720 10996 19748 11036
rect 21542 11024 21548 11076
rect 21600 11064 21606 11076
rect 22189 11067 22247 11073
rect 21600 11036 22140 11064
rect 21600 11024 21606 11036
rect 20622 10996 20628 11008
rect 19306 10968 19748 10996
rect 20583 10968 20628 10996
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 22112 10996 22140 11036
rect 22189 11033 22201 11067
rect 22235 11064 22247 11067
rect 22278 11064 22284 11076
rect 22235 11036 22284 11064
rect 22235 11033 22247 11036
rect 22189 11027 22247 11033
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 22405 11067 22463 11073
rect 22405 11064 22417 11067
rect 22388 11033 22417 11064
rect 22451 11064 22463 11067
rect 22756 11064 22784 11104
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23382 11141 23388 11144
rect 23201 11135 23259 11141
rect 23201 11132 23213 11135
rect 23072 11104 23213 11132
rect 23072 11092 23078 11104
rect 23201 11101 23213 11104
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23349 11135 23388 11141
rect 23349 11101 23361 11135
rect 23349 11095 23388 11101
rect 23382 11092 23388 11095
rect 23440 11092 23446 11144
rect 23707 11135 23765 11141
rect 23707 11101 23719 11135
rect 23753 11132 23765 11135
rect 24486 11132 24492 11144
rect 23753 11104 24348 11132
rect 24447 11104 24492 11132
rect 23753 11101 23765 11104
rect 23707 11095 23765 11101
rect 23477 11067 23535 11073
rect 23477 11064 23489 11067
rect 22451 11036 22692 11064
rect 22756 11036 23489 11064
rect 22451 11033 22463 11036
rect 22388 11027 22463 11033
rect 22388 10996 22416 11027
rect 22112 10968 22416 10996
rect 22664 10996 22692 11036
rect 23477 11033 23489 11036
rect 23523 11033 23535 11067
rect 23477 11027 23535 11033
rect 23569 11067 23627 11073
rect 23569 11033 23581 11067
rect 23615 11033 23627 11067
rect 24320 11064 24348 11104
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 24596 11141 24624 11172
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11132 24823 11135
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 24811 11104 25605 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 25593 11101 25605 11104
rect 25639 11101 25651 11135
rect 26326 11132 26332 11144
rect 26287 11104 26332 11132
rect 25593 11095 25651 11101
rect 26326 11092 26332 11104
rect 26384 11092 26390 11144
rect 26436 11132 26464 11172
rect 30190 11160 30196 11212
rect 30248 11200 30254 11212
rect 31113 11203 31171 11209
rect 31113 11200 31125 11203
rect 30248 11172 31125 11200
rect 30248 11160 30254 11172
rect 31113 11169 31125 11172
rect 31159 11169 31171 11203
rect 33428 11200 33456 11231
rect 31113 11163 31171 11169
rect 32600 11172 33456 11200
rect 26585 11135 26643 11141
rect 26585 11132 26597 11135
rect 26436 11104 26597 11132
rect 26585 11101 26597 11104
rect 26631 11101 26643 11135
rect 26585 11095 26643 11101
rect 31380 11135 31438 11141
rect 31380 11101 31392 11135
rect 31426 11132 31438 11135
rect 32600 11132 32628 11172
rect 32950 11132 32956 11144
rect 31426 11104 32628 11132
rect 32911 11104 32956 11132
rect 31426 11101 31438 11104
rect 31380 11095 31438 11101
rect 32950 11092 32956 11104
rect 33008 11092 33014 11144
rect 33318 11092 33324 11144
rect 33376 11132 33382 11144
rect 33413 11135 33471 11141
rect 33413 11132 33425 11135
rect 33376 11104 33425 11132
rect 33376 11092 33382 11104
rect 33413 11101 33425 11104
rect 33459 11101 33471 11135
rect 33413 11095 33471 11101
rect 25774 11064 25780 11076
rect 24320 11036 25780 11064
rect 23569 11027 23627 11033
rect 23290 10996 23296 11008
rect 22664 10968 23296 10996
rect 23290 10956 23296 10968
rect 23348 10956 23354 11008
rect 23584 10996 23612 11027
rect 25774 11024 25780 11036
rect 25832 11024 25838 11076
rect 32122 11024 32128 11076
rect 32180 11064 32186 11076
rect 33520 11064 33548 11240
rect 43254 11228 43260 11240
rect 43312 11228 43318 11280
rect 35621 11203 35679 11209
rect 35621 11169 35633 11203
rect 35667 11200 35679 11203
rect 37550 11200 37556 11212
rect 35667 11172 37556 11200
rect 35667 11169 35679 11172
rect 35621 11163 35679 11169
rect 37550 11160 37556 11172
rect 37608 11160 37614 11212
rect 40862 11160 40868 11212
rect 40920 11200 40926 11212
rect 40957 11203 41015 11209
rect 40957 11200 40969 11203
rect 40920 11172 40969 11200
rect 40920 11160 40926 11172
rect 40957 11169 40969 11172
rect 41003 11169 41015 11203
rect 40957 11163 41015 11169
rect 47780 11157 47808 11308
rect 48590 11296 48596 11308
rect 48648 11296 48654 11348
rect 50890 11336 50896 11348
rect 50851 11308 50896 11336
rect 50890 11296 50896 11308
rect 50948 11296 50954 11348
rect 51077 11339 51135 11345
rect 51077 11305 51089 11339
rect 51123 11336 51135 11339
rect 51534 11336 51540 11348
rect 51123 11308 51540 11336
rect 51123 11305 51135 11308
rect 51077 11299 51135 11305
rect 51534 11296 51540 11308
rect 51592 11296 51598 11348
rect 47765 11151 47823 11157
rect 35345 11135 35403 11141
rect 35345 11101 35357 11135
rect 35391 11132 35403 11135
rect 35710 11132 35716 11144
rect 35391 11104 35716 11132
rect 35391 11101 35403 11104
rect 35345 11095 35403 11101
rect 35710 11092 35716 11104
rect 35768 11092 35774 11144
rect 36262 11132 36268 11144
rect 36223 11104 36268 11132
rect 36262 11092 36268 11104
rect 36320 11092 36326 11144
rect 36354 11092 36360 11144
rect 36412 11132 36418 11144
rect 36538 11132 36544 11144
rect 36412 11104 36457 11132
rect 36499 11104 36544 11132
rect 36412 11092 36418 11104
rect 36538 11092 36544 11104
rect 36596 11092 36602 11144
rect 36633 11135 36691 11141
rect 36633 11101 36645 11135
rect 36679 11132 36691 11135
rect 38470 11132 38476 11144
rect 36679 11104 38476 11132
rect 36679 11101 36691 11104
rect 36633 11095 36691 11101
rect 38470 11092 38476 11104
rect 38528 11092 38534 11144
rect 41141 11135 41199 11141
rect 41141 11101 41153 11135
rect 41187 11132 41199 11135
rect 41506 11132 41512 11144
rect 41187 11104 41512 11132
rect 41187 11101 41199 11104
rect 41141 11095 41199 11101
rect 41506 11092 41512 11104
rect 41564 11132 41570 11144
rect 43714 11132 43720 11144
rect 41564 11104 43720 11132
rect 41564 11092 41570 11104
rect 43714 11092 43720 11104
rect 43772 11092 43778 11144
rect 47765 11117 47777 11151
rect 47811 11117 47823 11151
rect 47765 11111 47823 11117
rect 48225 11135 48283 11141
rect 48225 11101 48237 11135
rect 48271 11101 48283 11135
rect 48481 11135 48539 11141
rect 48481 11132 48493 11135
rect 48225 11095 48283 11101
rect 48424 11104 48493 11132
rect 41325 11067 41383 11073
rect 41325 11064 41337 11067
rect 32180 11036 33548 11064
rect 38626 11036 41337 11064
rect 32180 11024 32186 11036
rect 23658 10996 23664 11008
rect 23584 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 28442 10956 28448 11008
rect 28500 10996 28506 11008
rect 28902 10996 28908 11008
rect 28500 10968 28908 10996
rect 28500 10956 28506 10968
rect 28902 10956 28908 10968
rect 28960 10956 28966 11008
rect 33042 10996 33048 11008
rect 33003 10968 33048 10996
rect 33042 10956 33048 10968
rect 33100 10956 33106 11008
rect 33137 10999 33195 11005
rect 33137 10965 33149 10999
rect 33183 10996 33195 10999
rect 33226 10996 33232 11008
rect 33183 10968 33232 10996
rect 33183 10965 33195 10968
rect 33137 10959 33195 10965
rect 33226 10956 33232 10968
rect 33284 10956 33290 11008
rect 36078 10996 36084 11008
rect 36039 10968 36084 10996
rect 36078 10956 36084 10968
rect 36136 10956 36142 11008
rect 36354 10956 36360 11008
rect 36412 10996 36418 11008
rect 38626 10996 38654 11036
rect 41325 11033 41337 11036
rect 41371 11033 41383 11067
rect 41325 11027 41383 11033
rect 42426 11024 42432 11076
rect 42484 11064 42490 11076
rect 42484 11036 42932 11064
rect 42484 11024 42490 11036
rect 36412 10968 38654 10996
rect 42904 10996 42932 11036
rect 45554 11024 45560 11076
rect 45612 11064 45618 11076
rect 48240 11064 48268 11095
rect 48314 11064 48320 11076
rect 45612 11036 48320 11064
rect 45612 11024 45618 11036
rect 48314 11024 48320 11036
rect 48372 11024 48378 11076
rect 42978 10996 42984 11008
rect 42904 10968 42984 10996
rect 36412 10956 36418 10968
rect 42978 10956 42984 10968
rect 43036 10956 43042 11008
rect 47581 10999 47639 11005
rect 47581 10965 47593 10999
rect 47627 10996 47639 10999
rect 48424 10996 48452 11104
rect 48481 11101 48493 11104
rect 48527 11101 48539 11135
rect 53469 11135 53527 11141
rect 53469 11132 53481 11135
rect 48481 11095 48539 11101
rect 51046 11104 53481 11132
rect 50709 11067 50767 11073
rect 50709 11033 50721 11067
rect 50755 11064 50767 11067
rect 51046 11064 51074 11104
rect 53469 11101 53481 11104
rect 53515 11132 53527 11135
rect 54386 11132 54392 11144
rect 53515 11104 54392 11132
rect 53515 11101 53527 11104
rect 53469 11095 53527 11101
rect 54386 11092 54392 11104
rect 54444 11092 54450 11144
rect 50755 11036 51074 11064
rect 50755 11033 50767 11036
rect 50709 11027 50767 11033
rect 47627 10968 48452 10996
rect 49605 10999 49663 11005
rect 47627 10965 47639 10968
rect 47581 10959 47639 10965
rect 49605 10965 49617 10999
rect 49651 10996 49663 10999
rect 49878 10996 49884 11008
rect 49651 10968 49884 10996
rect 49651 10965 49663 10968
rect 49605 10959 49663 10965
rect 49878 10956 49884 10968
rect 49936 10996 49942 11008
rect 50909 10999 50967 11005
rect 50909 10996 50921 10999
rect 49936 10968 50921 10996
rect 49936 10956 49942 10968
rect 50909 10965 50921 10968
rect 50955 10965 50967 10999
rect 50909 10959 50967 10965
rect 53098 10956 53104 11008
rect 53156 10996 53162 11008
rect 53561 10999 53619 11005
rect 53561 10996 53573 10999
rect 53156 10968 53573 10996
rect 53156 10956 53162 10968
rect 53561 10965 53573 10968
rect 53607 10965 53619 10999
rect 53561 10959 53619 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 6917 10795 6975 10801
rect 6917 10761 6929 10795
rect 6963 10792 6975 10795
rect 7006 10792 7012 10804
rect 6963 10764 7012 10792
rect 6963 10761 6975 10764
rect 6917 10755 6975 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11112 10764 22094 10792
rect 11112 10752 11118 10764
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3568 10696 9352 10724
rect 3568 10684 3574 10696
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2314 10665 2320 10668
rect 2308 10656 2320 10665
rect 2275 10628 2320 10656
rect 2308 10619 2320 10628
rect 2314 10616 2320 10619
rect 2372 10616 2378 10668
rect 7098 10656 7104 10668
rect 7011 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7374 10656 7380 10668
rect 7335 10628 7380 10656
rect 7374 10616 7380 10628
rect 7432 10616 7438 10668
rect 6914 10588 6920 10600
rect 6886 10548 6920 10588
rect 6972 10548 6978 10600
rect 3602 10520 3608 10532
rect 3252 10492 3608 10520
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 3252 10452 3280 10492
rect 3602 10480 3608 10492
rect 3660 10480 3666 10532
rect 3418 10452 3424 10464
rect 1443 10424 3280 10452
rect 3331 10424 3424 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 3418 10412 3424 10424
rect 3476 10452 3482 10464
rect 6886 10452 6914 10548
rect 3476 10424 6914 10452
rect 7116 10452 7144 10616
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10588 7343 10591
rect 7484 10588 7512 10696
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7331 10560 7512 10588
rect 7576 10588 7604 10619
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 7892 10628 8125 10656
rect 7892 10616 7898 10628
rect 8113 10625 8125 10628
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 7742 10588 7748 10600
rect 7576 10560 7748 10588
rect 7331 10557 7343 10560
rect 7285 10551 7343 10557
rect 7742 10548 7748 10560
rect 7800 10588 7806 10600
rect 8297 10591 8355 10597
rect 8297 10588 8309 10591
rect 7800 10560 8309 10588
rect 7800 10548 7806 10560
rect 8297 10557 8309 10560
rect 8343 10557 8355 10591
rect 9324 10588 9352 10696
rect 10502 10684 10508 10736
rect 10560 10724 10566 10736
rect 10962 10724 10968 10736
rect 10560 10696 10968 10724
rect 10560 10684 10566 10696
rect 10962 10684 10968 10696
rect 11020 10724 11026 10736
rect 12069 10727 12127 10733
rect 11020 10696 11928 10724
rect 11020 10684 11026 10696
rect 11606 10656 11612 10668
rect 11567 10628 11612 10656
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 11698 10616 11704 10668
rect 11756 10656 11762 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11756 10628 11805 10656
rect 11756 10616 11762 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11900 10656 11928 10696
rect 12069 10693 12081 10727
rect 12115 10724 12127 10727
rect 14090 10724 14096 10736
rect 12115 10696 14096 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 14090 10684 14096 10696
rect 14148 10724 14154 10736
rect 14366 10724 14372 10736
rect 14148 10696 14372 10724
rect 14148 10684 14154 10696
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 14544 10727 14602 10733
rect 14544 10693 14556 10727
rect 14590 10724 14602 10727
rect 15010 10724 15016 10736
rect 14590 10696 15016 10724
rect 14590 10693 14602 10696
rect 14544 10687 14602 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 16390 10724 16396 10736
rect 15252 10696 16396 10724
rect 15252 10684 15258 10696
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17313 10727 17371 10733
rect 17313 10693 17325 10727
rect 17359 10724 17371 10727
rect 17678 10724 17684 10736
rect 17359 10696 17684 10724
rect 17359 10693 17371 10696
rect 17313 10687 17371 10693
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 19153 10727 19211 10733
rect 19153 10693 19165 10727
rect 19199 10724 19211 10727
rect 19426 10724 19432 10736
rect 19199 10696 19432 10724
rect 19199 10693 19211 10696
rect 19153 10687 19211 10693
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 19518 10684 19524 10736
rect 19576 10724 19582 10736
rect 20622 10724 20628 10736
rect 19576 10696 20628 10724
rect 19576 10684 19582 10696
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 22066 10724 22094 10764
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 23382 10792 23388 10804
rect 22428 10764 23388 10792
rect 22428 10752 22434 10764
rect 23382 10752 23388 10764
rect 23440 10792 23446 10804
rect 27338 10792 27344 10804
rect 23440 10764 27344 10792
rect 23440 10752 23446 10764
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 31481 10795 31539 10801
rect 31481 10761 31493 10795
rect 31527 10792 31539 10795
rect 33042 10792 33048 10804
rect 31527 10764 33048 10792
rect 31527 10761 31539 10764
rect 31481 10755 31539 10761
rect 33042 10752 33048 10764
rect 33100 10752 33106 10804
rect 38746 10752 38752 10804
rect 38804 10792 38810 10804
rect 41966 10792 41972 10804
rect 38804 10764 41972 10792
rect 38804 10752 38810 10764
rect 41966 10752 41972 10764
rect 42024 10792 42030 10804
rect 44542 10792 44548 10804
rect 42024 10764 44548 10792
rect 42024 10752 42030 10764
rect 44542 10752 44548 10764
rect 44600 10752 44606 10804
rect 48498 10752 48504 10804
rect 48556 10792 48562 10804
rect 48869 10795 48927 10801
rect 48869 10792 48881 10795
rect 48556 10764 48881 10792
rect 48556 10752 48562 10764
rect 48869 10761 48881 10764
rect 48915 10761 48927 10795
rect 48869 10755 48927 10761
rect 50249 10795 50307 10801
rect 50249 10761 50261 10795
rect 50295 10792 50307 10795
rect 50798 10792 50804 10804
rect 50295 10764 50804 10792
rect 50295 10761 50307 10764
rect 50249 10755 50307 10761
rect 50798 10752 50804 10764
rect 50856 10752 50862 10804
rect 54386 10792 54392 10804
rect 54347 10764 54392 10792
rect 54386 10752 54392 10764
rect 54444 10752 54450 10804
rect 35526 10724 35532 10736
rect 22066 10696 35532 10724
rect 35526 10684 35532 10696
rect 35584 10684 35590 10736
rect 48590 10724 48596 10736
rect 36556 10696 48596 10724
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 11900 10628 12357 10656
rect 11793 10619 11851 10625
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 14274 10656 14280 10668
rect 14235 10628 14280 10656
rect 12345 10619 12403 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 17126 10656 17132 10668
rect 16632 10628 17132 10656
rect 16632 10616 16638 10628
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 19337 10659 19395 10665
rect 19337 10625 19349 10659
rect 19383 10656 19395 10659
rect 19613 10659 19671 10665
rect 19383 10628 19564 10656
rect 19383 10625 19395 10628
rect 19337 10619 19395 10625
rect 19536 10600 19564 10628
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19613 10619 19671 10625
rect 13998 10588 14004 10600
rect 9324 10560 14004 10588
rect 8297 10551 8355 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 19518 10548 19524 10600
rect 19576 10548 19582 10600
rect 7193 10523 7251 10529
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 7926 10520 7932 10532
rect 7239 10492 7932 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 7760 10464 7788 10492
rect 7926 10480 7932 10492
rect 7984 10480 7990 10532
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 10870 10520 10876 10532
rect 10560 10492 10876 10520
rect 10560 10480 10566 10492
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 16390 10480 16396 10532
rect 16448 10520 16454 10532
rect 19150 10520 19156 10532
rect 16448 10492 19156 10520
rect 16448 10480 16454 10492
rect 19150 10480 19156 10492
rect 19208 10520 19214 10532
rect 19628 10520 19656 10619
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 30929 10659 30987 10665
rect 30929 10656 30941 10659
rect 27672 10628 30941 10656
rect 27672 10616 27678 10628
rect 30929 10625 30941 10628
rect 30975 10625 30987 10659
rect 30929 10619 30987 10625
rect 31297 10659 31355 10665
rect 31297 10625 31309 10659
rect 31343 10656 31355 10659
rect 32122 10656 32128 10668
rect 31343 10628 32128 10656
rect 31343 10625 31355 10628
rect 31297 10619 31355 10625
rect 32122 10616 32128 10628
rect 32180 10616 32186 10668
rect 36078 10656 36084 10668
rect 36039 10628 36084 10656
rect 36078 10616 36084 10628
rect 36136 10616 36142 10668
rect 36354 10656 36360 10668
rect 36315 10628 36360 10656
rect 36354 10616 36360 10628
rect 36412 10616 36418 10668
rect 36556 10665 36584 10696
rect 48590 10684 48596 10696
rect 48648 10724 48654 10736
rect 49878 10724 49884 10736
rect 48648 10696 49280 10724
rect 49839 10696 49884 10724
rect 48648 10684 48654 10696
rect 36541 10659 36599 10665
rect 36541 10625 36553 10659
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 30190 10548 30196 10600
rect 30248 10588 30254 10600
rect 36556 10588 36584 10619
rect 42334 10616 42340 10668
rect 42392 10656 42398 10668
rect 49252 10665 49280 10696
rect 49878 10684 49884 10696
rect 49936 10684 49942 10736
rect 49970 10684 49976 10736
rect 50028 10724 50034 10736
rect 50081 10727 50139 10733
rect 50081 10724 50093 10727
rect 50028 10696 50093 10724
rect 50028 10684 50034 10696
rect 50081 10693 50093 10696
rect 50127 10693 50139 10727
rect 50081 10687 50139 10693
rect 42889 10659 42947 10665
rect 42889 10656 42901 10659
rect 42392 10628 42901 10656
rect 42392 10616 42398 10628
rect 42889 10625 42901 10628
rect 42935 10625 42947 10659
rect 42889 10619 42947 10625
rect 49237 10659 49295 10665
rect 49237 10625 49249 10659
rect 49283 10625 49295 10659
rect 49237 10619 49295 10625
rect 49329 10659 49387 10665
rect 49329 10625 49341 10659
rect 49375 10656 49387 10659
rect 49896 10656 49924 10684
rect 53282 10665 53288 10668
rect 49375 10628 49924 10656
rect 49375 10625 49387 10628
rect 49329 10619 49387 10625
rect 53276 10619 53288 10665
rect 53340 10656 53346 10668
rect 53340 10628 53376 10656
rect 53282 10616 53288 10619
rect 53340 10616 53346 10628
rect 30248 10560 36584 10588
rect 30248 10548 30254 10560
rect 48222 10548 48228 10600
rect 48280 10588 48286 10600
rect 49053 10591 49111 10597
rect 49053 10588 49065 10591
rect 48280 10560 49065 10588
rect 48280 10548 48286 10560
rect 49053 10557 49065 10560
rect 49099 10557 49111 10591
rect 49053 10551 49111 10557
rect 49145 10591 49203 10597
rect 49145 10557 49157 10591
rect 49191 10588 49203 10591
rect 49191 10560 50108 10588
rect 49191 10557 49203 10560
rect 49145 10551 49203 10557
rect 19208 10492 19656 10520
rect 31312 10492 31524 10520
rect 19208 10480 19214 10492
rect 7558 10452 7564 10464
rect 7116 10424 7564 10452
rect 3476 10412 3482 10424
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 7742 10412 7748 10464
rect 7800 10412 7806 10464
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 11664 10424 15669 10452
rect 11664 10412 11670 10424
rect 15657 10421 15669 10424
rect 15703 10452 15715 10455
rect 16022 10452 16028 10464
rect 15703 10424 16028 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 31312 10461 31340 10492
rect 31297 10455 31355 10461
rect 31297 10421 31309 10455
rect 31343 10421 31355 10455
rect 31496 10452 31524 10492
rect 31570 10480 31576 10532
rect 31628 10520 31634 10532
rect 33410 10520 33416 10532
rect 31628 10492 33416 10520
rect 31628 10480 31634 10492
rect 33410 10480 33416 10492
rect 33468 10480 33474 10532
rect 50080 10464 50108 10560
rect 52638 10548 52644 10600
rect 52696 10588 52702 10600
rect 53009 10591 53067 10597
rect 53009 10588 53021 10591
rect 52696 10560 53021 10588
rect 52696 10548 52702 10560
rect 53009 10557 53021 10560
rect 53055 10557 53067 10591
rect 53009 10551 53067 10557
rect 32214 10452 32220 10464
rect 31496 10424 32220 10452
rect 31297 10415 31355 10421
rect 32214 10412 32220 10424
rect 32272 10412 32278 10464
rect 35894 10452 35900 10464
rect 35855 10424 35900 10452
rect 35894 10412 35900 10424
rect 35952 10412 35958 10464
rect 42705 10455 42763 10461
rect 42705 10421 42717 10455
rect 42751 10452 42763 10455
rect 43070 10452 43076 10464
rect 42751 10424 43076 10452
rect 42751 10421 42763 10424
rect 42705 10415 42763 10421
rect 43070 10412 43076 10424
rect 43128 10412 43134 10464
rect 50062 10452 50068 10464
rect 49975 10424 50068 10452
rect 50062 10412 50068 10424
rect 50120 10452 50126 10464
rect 50982 10452 50988 10464
rect 50120 10424 50988 10452
rect 50120 10412 50126 10424
rect 50982 10412 50988 10424
rect 51040 10412 51046 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2406 10248 2412 10260
rect 2271 10220 2412 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 6144 10220 6193 10248
rect 6144 10208 6150 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 11698 10208 11704 10260
rect 11756 10248 11762 10260
rect 11974 10248 11980 10260
rect 11756 10220 11980 10248
rect 11756 10208 11762 10220
rect 11974 10208 11980 10220
rect 12032 10248 12038 10260
rect 12032 10220 12204 10248
rect 12032 10208 12038 10220
rect 2590 10140 2596 10192
rect 2648 10140 2654 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 10192 10152 12081 10180
rect 10192 10140 10198 10152
rect 12069 10149 12081 10152
rect 12115 10149 12127 10183
rect 12176 10180 12204 10220
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14642 10248 14648 10260
rect 14332 10220 14648 10248
rect 14332 10208 14338 10220
rect 14642 10208 14648 10220
rect 14700 10248 14706 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14700 10220 15025 10248
rect 14700 10208 14706 10220
rect 15013 10217 15025 10220
rect 15059 10248 15071 10251
rect 15059 10220 16712 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15197 10183 15255 10189
rect 15197 10180 15209 10183
rect 12176 10152 15209 10180
rect 12069 10143 12127 10149
rect 15197 10149 15209 10152
rect 15243 10149 15255 10183
rect 15197 10143 15255 10149
rect 2608 10112 2636 10140
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2608 10084 2789 10112
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 4801 10115 4859 10121
rect 4801 10112 4813 10115
rect 3844 10084 4813 10112
rect 3844 10072 3850 10084
rect 4801 10081 4813 10084
rect 4847 10081 4859 10115
rect 4801 10075 4859 10081
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7834 10112 7840 10124
rect 7147 10084 7840 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 16574 10112 16580 10124
rect 11440 10084 16580 10112
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 3418 10044 3424 10056
rect 2639 10016 3424 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 4948 10016 6929 10044
rect 4948 10004 4954 10016
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 11440 10053 11468 10084
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 11606 10053 11612 10056
rect 11425 10047 11483 10053
rect 7248 10016 7293 10044
rect 7248 10004 7254 10016
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11573 10047 11612 10053
rect 11573 10013 11585 10047
rect 11573 10007 11612 10013
rect 11606 10004 11612 10007
rect 11664 10004 11670 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11756 10016 11801 10044
rect 11756 10004 11762 10016
rect 11882 10004 11888 10056
rect 11940 10053 11946 10056
rect 11940 10044 11948 10053
rect 11940 10016 11985 10044
rect 11940 10007 11948 10016
rect 11940 10004 11946 10007
rect 5068 9979 5126 9985
rect 5068 9945 5080 9979
rect 5114 9976 5126 9979
rect 6362 9976 6368 9988
rect 5114 9948 6368 9976
rect 5114 9945 5126 9948
rect 5068 9939 5126 9945
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9945 11851 9979
rect 14826 9976 14832 9988
rect 14787 9948 14832 9976
rect 11793 9939 11851 9945
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 2740 9880 2785 9908
rect 2740 9868 2746 9880
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6512 9880 6745 9908
rect 6512 9868 6518 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 11808 9908 11836 9939
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15045 9979 15103 9985
rect 15045 9945 15057 9979
rect 15091 9976 15103 9979
rect 15194 9976 15200 9988
rect 15091 9948 15200 9976
rect 15091 9945 15103 9948
rect 15045 9939 15103 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 16684 9976 16712 10220
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18141 10251 18199 10257
rect 18141 10248 18153 10251
rect 18104 10220 18153 10248
rect 18104 10208 18110 10220
rect 18141 10217 18153 10220
rect 18187 10217 18199 10251
rect 18141 10211 18199 10217
rect 34790 10208 34796 10260
rect 34848 10248 34854 10260
rect 34885 10251 34943 10257
rect 34885 10248 34897 10251
rect 34848 10220 34897 10248
rect 34848 10208 34854 10220
rect 34885 10217 34897 10220
rect 34931 10217 34943 10251
rect 36078 10248 36084 10260
rect 36039 10220 36084 10248
rect 34885 10211 34943 10217
rect 36078 10208 36084 10220
rect 36136 10248 36142 10260
rect 36722 10248 36728 10260
rect 36136 10220 36728 10248
rect 36136 10208 36142 10220
rect 36722 10208 36728 10220
rect 36780 10208 36786 10260
rect 42334 10248 42340 10260
rect 42295 10220 42340 10248
rect 42334 10208 42340 10220
rect 42392 10208 42398 10260
rect 47670 10248 47676 10260
rect 47631 10220 47676 10248
rect 47670 10208 47676 10220
rect 47728 10248 47734 10260
rect 49602 10248 49608 10260
rect 47728 10220 49608 10248
rect 47728 10208 47734 10220
rect 49602 10208 49608 10220
rect 49660 10208 49666 10260
rect 53282 10248 53288 10260
rect 53243 10220 53288 10248
rect 53282 10208 53288 10220
rect 53340 10208 53346 10260
rect 26878 10140 26884 10192
rect 26936 10180 26942 10192
rect 26936 10152 41276 10180
rect 26936 10140 26942 10152
rect 31938 10072 31944 10124
rect 31996 10112 32002 10124
rect 36538 10112 36544 10124
rect 31996 10084 32444 10112
rect 31996 10072 32002 10084
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 18230 10044 18236 10056
rect 17359 10016 18236 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 21174 10044 21180 10056
rect 19576 10016 21180 10044
rect 19576 10004 19582 10016
rect 21174 10004 21180 10016
rect 21232 10044 21238 10056
rect 26053 10047 26111 10053
rect 26053 10044 26065 10047
rect 21232 10016 26065 10044
rect 21232 10004 21238 10016
rect 26053 10013 26065 10016
rect 26099 10013 26111 10047
rect 26326 10044 26332 10056
rect 26287 10016 26332 10044
rect 26053 10007 26111 10013
rect 18049 9979 18107 9985
rect 18049 9976 18061 9979
rect 16684 9948 18061 9976
rect 18049 9945 18061 9948
rect 18095 9945 18107 9979
rect 26068 9976 26096 10007
rect 26326 10004 26332 10016
rect 26384 10004 26390 10056
rect 32416 10053 32444 10084
rect 34716 10084 36544 10112
rect 34716 10056 34744 10084
rect 36538 10072 36544 10084
rect 36596 10072 36602 10124
rect 32125 10047 32183 10053
rect 32125 10013 32137 10047
rect 32171 10013 32183 10047
rect 32125 10007 32183 10013
rect 32401 10047 32459 10053
rect 32401 10013 32413 10047
rect 32447 10013 32459 10047
rect 32401 10007 32459 10013
rect 32493 10047 32551 10053
rect 32493 10013 32505 10047
rect 32539 10044 32551 10047
rect 33502 10044 33508 10056
rect 32539 10016 33508 10044
rect 32539 10013 32551 10016
rect 32493 10007 32551 10013
rect 32030 9976 32036 9988
rect 26068 9948 32036 9976
rect 18049 9939 18107 9945
rect 32030 9936 32036 9948
rect 32088 9936 32094 9988
rect 10928 9880 11836 9908
rect 10928 9868 10934 9880
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17276 9880 17417 9908
rect 17276 9868 17282 9880
rect 17405 9877 17417 9880
rect 17451 9908 17463 9911
rect 18414 9908 18420 9920
rect 17451 9880 18420 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 25866 9908 25872 9920
rect 25827 9880 25872 9908
rect 25866 9868 25872 9880
rect 25924 9868 25930 9920
rect 26237 9911 26295 9917
rect 26237 9877 26249 9911
rect 26283 9908 26295 9911
rect 27062 9908 27068 9920
rect 26283 9880 27068 9908
rect 26283 9877 26295 9880
rect 26237 9871 26295 9877
rect 27062 9868 27068 9880
rect 27120 9908 27126 9920
rect 31570 9908 31576 9920
rect 27120 9880 31576 9908
rect 27120 9868 27126 9880
rect 31570 9868 31576 9880
rect 31628 9868 31634 9920
rect 32140 9908 32168 10007
rect 33502 10004 33508 10016
rect 33560 10004 33566 10056
rect 34698 10044 34704 10056
rect 34659 10016 34704 10044
rect 34698 10004 34704 10016
rect 34756 10004 34762 10056
rect 35713 10047 35771 10053
rect 35713 10013 35725 10047
rect 35759 10044 35771 10047
rect 37458 10044 37464 10056
rect 35759 10016 37464 10044
rect 35759 10013 35771 10016
rect 35713 10007 35771 10013
rect 37458 10004 37464 10016
rect 37516 10004 37522 10056
rect 38565 10047 38623 10053
rect 38565 10013 38577 10047
rect 38611 10044 38623 10047
rect 39206 10044 39212 10056
rect 38611 10016 39212 10044
rect 38611 10013 38623 10016
rect 38565 10007 38623 10013
rect 39206 10004 39212 10016
rect 39264 10004 39270 10056
rect 40954 10044 40960 10056
rect 40915 10016 40960 10044
rect 40954 10004 40960 10016
rect 41012 10004 41018 10056
rect 41248 10053 41276 10152
rect 42978 10112 42984 10124
rect 42939 10084 42984 10112
rect 42978 10072 42984 10084
rect 43036 10072 43042 10124
rect 45554 10072 45560 10124
rect 45612 10112 45618 10124
rect 45649 10115 45707 10121
rect 45649 10112 45661 10115
rect 45612 10084 45661 10112
rect 45612 10072 45618 10084
rect 45649 10081 45661 10084
rect 45695 10081 45707 10115
rect 45649 10075 45707 10081
rect 52914 10072 52920 10124
rect 52972 10112 52978 10124
rect 53285 10115 53343 10121
rect 53285 10112 53297 10115
rect 52972 10084 53297 10112
rect 52972 10072 52978 10084
rect 53285 10081 53297 10084
rect 53331 10081 53343 10115
rect 53285 10075 53343 10081
rect 41233 10047 41291 10053
rect 41233 10013 41245 10047
rect 41279 10013 41291 10047
rect 41233 10007 41291 10013
rect 41322 10004 41328 10056
rect 41380 10044 41386 10056
rect 41966 10044 41972 10056
rect 41380 10016 41425 10044
rect 41927 10016 41972 10044
rect 41380 10004 41386 10016
rect 41966 10004 41972 10016
rect 42024 10004 42030 10056
rect 42150 10044 42156 10056
rect 42111 10016 42156 10044
rect 42150 10004 42156 10016
rect 42208 10004 42214 10056
rect 43070 10004 43076 10056
rect 43128 10044 43134 10056
rect 43237 10047 43295 10053
rect 43237 10044 43249 10047
rect 43128 10016 43249 10044
rect 43128 10004 43134 10016
rect 43237 10013 43249 10016
rect 43283 10013 43295 10047
rect 47581 10047 47639 10053
rect 47581 10044 47593 10047
rect 43237 10007 43295 10013
rect 47044 10016 47593 10044
rect 32306 9976 32312 9988
rect 32267 9948 32312 9976
rect 32306 9936 32312 9948
rect 32364 9936 32370 9988
rect 33134 9976 33140 9988
rect 32508 9948 33140 9976
rect 32508 9908 32536 9948
rect 33134 9936 33140 9948
rect 33192 9936 33198 9988
rect 36081 9979 36139 9985
rect 36081 9945 36093 9979
rect 36127 9976 36139 9979
rect 36170 9976 36176 9988
rect 36127 9948 36176 9976
rect 36127 9945 36139 9948
rect 36081 9939 36139 9945
rect 36170 9936 36176 9948
rect 36228 9936 36234 9988
rect 41141 9979 41199 9985
rect 41141 9945 41153 9979
rect 41187 9945 41199 9979
rect 41141 9939 41199 9945
rect 32674 9908 32680 9920
rect 32140 9880 32536 9908
rect 32635 9880 32680 9908
rect 32674 9868 32680 9880
rect 32732 9868 32738 9920
rect 35250 9868 35256 9920
rect 35308 9908 35314 9920
rect 35618 9908 35624 9920
rect 35308 9880 35624 9908
rect 35308 9868 35314 9880
rect 35618 9868 35624 9880
rect 35676 9868 35682 9920
rect 36262 9908 36268 9920
rect 36223 9880 36268 9908
rect 36262 9868 36268 9880
rect 36320 9868 36326 9920
rect 38010 9868 38016 9920
rect 38068 9908 38074 9920
rect 38381 9911 38439 9917
rect 38381 9908 38393 9911
rect 38068 9880 38393 9908
rect 38068 9868 38074 9880
rect 38381 9877 38393 9880
rect 38427 9877 38439 9911
rect 41156 9908 41184 9939
rect 45554 9936 45560 9988
rect 45612 9976 45618 9988
rect 45894 9979 45952 9985
rect 45894 9976 45906 9979
rect 45612 9948 45906 9976
rect 45612 9936 45618 9948
rect 45894 9945 45906 9948
rect 45940 9945 45952 9979
rect 45894 9939 45952 9945
rect 47044 9920 47072 10016
rect 47581 10013 47593 10016
rect 47627 10013 47639 10047
rect 53098 10044 53104 10056
rect 53059 10016 53104 10044
rect 47581 10007 47639 10013
rect 53098 10004 53104 10016
rect 53156 10004 53162 10056
rect 53190 10004 53196 10056
rect 53248 10044 53254 10056
rect 53248 10016 53293 10044
rect 53248 10004 53254 10016
rect 52917 9979 52975 9985
rect 52917 9945 52929 9979
rect 52963 9976 52975 9979
rect 53926 9976 53932 9988
rect 52963 9948 53932 9976
rect 52963 9945 52975 9948
rect 52917 9939 52975 9945
rect 53926 9936 53932 9948
rect 53984 9936 53990 9988
rect 41414 9908 41420 9920
rect 41156 9880 41420 9908
rect 38381 9871 38439 9877
rect 41414 9868 41420 9880
rect 41472 9868 41478 9920
rect 41506 9868 41512 9920
rect 41564 9908 41570 9920
rect 41564 9880 41609 9908
rect 41564 9868 41570 9880
rect 43898 9868 43904 9920
rect 43956 9908 43962 9920
rect 44361 9911 44419 9917
rect 44361 9908 44373 9911
rect 43956 9880 44373 9908
rect 43956 9868 43962 9880
rect 44361 9877 44373 9880
rect 44407 9877 44419 9911
rect 47026 9908 47032 9920
rect 46987 9880 47032 9908
rect 44361 9871 44419 9877
rect 47026 9868 47032 9880
rect 47084 9868 47090 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6144 9676 6745 9704
rect 6144 9664 6150 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 11882 9704 11888 9716
rect 6733 9667 6791 9673
rect 8128 9676 11888 9704
rect 6362 9636 6368 9648
rect 6323 9608 6368 9636
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 8128 9645 8156 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 12342 9704 12348 9716
rect 12176 9676 12348 9704
rect 8113 9639 8171 9645
rect 8113 9605 8125 9639
rect 8159 9605 8171 9639
rect 10594 9636 10600 9648
rect 8113 9599 8171 9605
rect 9048 9608 10600 9636
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 3234 9568 3240 9580
rect 1443 9540 3240 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7466 9568 7472 9580
rect 6871 9540 7472 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 6564 9500 6592 9531
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 8846 9568 8852 9580
rect 8807 9540 8852 9568
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 9048 9577 9076 9608
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 12176 9645 12204 9676
rect 12342 9664 12348 9676
rect 12400 9704 12406 9716
rect 14826 9704 14832 9716
rect 12400 9676 14832 9704
rect 12400 9664 12406 9676
rect 14826 9664 14832 9676
rect 14884 9704 14890 9716
rect 18230 9704 18236 9716
rect 14884 9676 18236 9704
rect 14884 9664 14890 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 32030 9664 32036 9716
rect 32088 9704 32094 9716
rect 38654 9704 38660 9716
rect 32088 9676 38660 9704
rect 32088 9664 32094 9676
rect 38654 9664 38660 9676
rect 38712 9664 38718 9716
rect 39206 9664 39212 9716
rect 39264 9704 39270 9716
rect 41509 9707 41567 9713
rect 39264 9676 39344 9704
rect 39264 9664 39270 9676
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11020 9608 11989 9636
rect 11020 9596 11026 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 12161 9639 12219 9645
rect 12161 9605 12173 9639
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 17126 9636 17132 9648
rect 14608 9608 17132 9636
rect 14608 9596 14614 9608
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 25216 9639 25274 9645
rect 17236 9608 25176 9636
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9858 9568 9864 9580
rect 9819 9540 9864 9568
rect 9033 9531 9091 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 10008 9540 13277 9568
rect 10008 9528 10014 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 13354 9528 13360 9580
rect 13412 9568 13418 9580
rect 14274 9568 14280 9580
rect 13412 9540 13457 9568
rect 14235 9540 14280 9568
rect 13412 9528 13418 9540
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 16666 9568 16672 9580
rect 16627 9540 16672 9568
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 11698 9500 11704 9512
rect 6564 9472 11704 9500
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 13044 9472 13093 9500
rect 13044 9460 13050 9472
rect 13081 9469 13093 9472
rect 13127 9500 13139 9503
rect 13906 9500 13912 9512
rect 13127 9472 13912 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 13906 9460 13912 9472
rect 13964 9460 13970 9512
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 14642 9500 14648 9512
rect 14599 9472 14648 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17034 9500 17040 9512
rect 16991 9472 17040 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 17236 9432 17264 9608
rect 18230 9568 18236 9580
rect 18191 9540 18236 9568
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9568 19303 9571
rect 19334 9568 19340 9580
rect 19291 9540 19340 9568
rect 19291 9537 19303 9540
rect 19245 9531 19303 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19512 9571 19570 9577
rect 19512 9537 19524 9571
rect 19558 9568 19570 9571
rect 20070 9568 20076 9580
rect 19558 9540 20076 9568
rect 19558 9537 19570 9540
rect 19512 9531 19570 9537
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 22370 9577 22376 9580
rect 22364 9531 22376 9577
rect 22428 9568 22434 9580
rect 25148 9568 25176 9608
rect 25216 9605 25228 9639
rect 25262 9636 25274 9639
rect 25866 9636 25872 9648
rect 25262 9608 25872 9636
rect 25262 9605 25274 9608
rect 25216 9599 25274 9605
rect 25866 9596 25872 9608
rect 25924 9596 25930 9648
rect 28436 9639 28494 9645
rect 28436 9605 28448 9639
rect 28482 9636 28494 9639
rect 32398 9636 32404 9648
rect 28482 9608 32404 9636
rect 28482 9605 28494 9608
rect 28436 9599 28494 9605
rect 32398 9596 32404 9608
rect 32456 9596 32462 9648
rect 39316 9645 39344 9676
rect 41509 9673 41521 9707
rect 41555 9704 41567 9707
rect 42150 9704 42156 9716
rect 41555 9676 42156 9704
rect 41555 9673 41567 9676
rect 41509 9667 41567 9673
rect 42150 9664 42156 9676
rect 42208 9664 42214 9716
rect 50706 9704 50712 9716
rect 50667 9676 50712 9704
rect 50706 9664 50712 9676
rect 50764 9664 50770 9716
rect 52638 9664 52644 9716
rect 52696 9704 52702 9716
rect 53558 9704 53564 9716
rect 52696 9676 53564 9704
rect 52696 9664 52702 9676
rect 53558 9664 53564 9676
rect 53616 9664 53622 9716
rect 56321 9707 56379 9713
rect 56321 9673 56333 9707
rect 56367 9673 56379 9707
rect 56321 9667 56379 9673
rect 33321 9639 33379 9645
rect 33321 9636 33333 9639
rect 33244 9608 33333 9636
rect 26878 9568 26884 9580
rect 22428 9540 22464 9568
rect 25148 9540 26884 9568
rect 22370 9528 22376 9531
rect 22428 9528 22434 9540
rect 26878 9528 26884 9540
rect 26936 9528 26942 9580
rect 29546 9528 29552 9580
rect 29604 9568 29610 9580
rect 30009 9571 30067 9577
rect 30009 9568 30021 9571
rect 29604 9540 30021 9568
rect 29604 9528 29610 9540
rect 30009 9537 30021 9540
rect 30055 9537 30067 9571
rect 30009 9531 30067 9537
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9568 31447 9571
rect 32674 9568 32680 9580
rect 31435 9540 32680 9568
rect 31435 9537 31447 9540
rect 31389 9531 31447 9537
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 33134 9568 33140 9580
rect 33095 9540 33140 9568
rect 33134 9528 33140 9540
rect 33192 9528 33198 9580
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18104 9472 18153 9500
rect 18104 9460 18110 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 17678 9432 17684 9444
rect 10652 9404 17264 9432
rect 17328 9404 17684 9432
rect 10652 9392 10658 9404
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 7524 9336 8217 9364
rect 7524 9324 7530 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8444 9336 8861 9364
rect 8444 9324 8450 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 8849 9327 8907 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10502 9364 10508 9376
rect 10008 9336 10508 9364
rect 10008 9324 10014 9336
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 13538 9364 13544 9376
rect 13499 9336 13544 9364
rect 13538 9324 13544 9336
rect 13596 9324 13602 9376
rect 14366 9324 14372 9376
rect 14424 9364 14430 9376
rect 16850 9364 16856 9376
rect 14424 9336 16856 9364
rect 14424 9324 14430 9336
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17328 9364 17356 9404
rect 17678 9392 17684 9404
rect 17736 9432 17742 9444
rect 18064 9432 18092 9460
rect 17736 9404 18092 9432
rect 17736 9392 17742 9404
rect 17000 9336 17356 9364
rect 17000 9324 17006 9336
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 17957 9367 18015 9373
rect 17957 9364 17969 9367
rect 17828 9336 17969 9364
rect 17828 9324 17834 9336
rect 17957 9333 17969 9336
rect 18003 9333 18015 9367
rect 18340 9364 18368 9463
rect 18414 9460 18420 9512
rect 18472 9500 18478 9512
rect 18472 9472 18517 9500
rect 18472 9460 18478 9472
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 22060 9472 22109 9500
rect 22060 9460 22066 9472
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 23474 9460 23480 9512
rect 23532 9500 23538 9512
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 23532 9472 24961 9500
rect 23532 9460 23538 9472
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 26786 9460 26792 9512
rect 26844 9500 26850 9512
rect 28166 9500 28172 9512
rect 26844 9472 28172 9500
rect 26844 9460 26850 9472
rect 28166 9460 28172 9472
rect 28224 9460 28230 9512
rect 31205 9503 31263 9509
rect 31205 9469 31217 9503
rect 31251 9500 31263 9503
rect 31754 9500 31760 9512
rect 31251 9472 31760 9500
rect 31251 9469 31263 9472
rect 31205 9463 31263 9469
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 26234 9392 26240 9444
rect 26292 9432 26298 9444
rect 26329 9435 26387 9441
rect 26329 9432 26341 9435
rect 26292 9404 26341 9432
rect 26292 9392 26298 9404
rect 26329 9401 26341 9404
rect 26375 9432 26387 9435
rect 27338 9432 27344 9444
rect 26375 9404 27344 9432
rect 26375 9401 26387 9404
rect 26329 9395 26387 9401
rect 27338 9392 27344 9404
rect 27396 9392 27402 9444
rect 33042 9392 33048 9444
rect 33100 9432 33106 9444
rect 33244 9432 33272 9608
rect 33321 9605 33333 9608
rect 33367 9605 33379 9639
rect 33321 9599 33379 9605
rect 38105 9639 38163 9645
rect 38105 9605 38117 9639
rect 38151 9605 38163 9639
rect 38105 9599 38163 9605
rect 39301 9639 39359 9645
rect 39301 9605 39313 9639
rect 39347 9605 39359 9639
rect 41230 9636 41236 9648
rect 41191 9608 41236 9636
rect 39301 9599 39359 9605
rect 33413 9571 33471 9577
rect 33413 9537 33425 9571
rect 33459 9537 33471 9571
rect 33413 9531 33471 9537
rect 33100 9404 33272 9432
rect 33100 9392 33106 9404
rect 20622 9364 20628 9376
rect 18340 9336 20628 9364
rect 17957 9327 18015 9333
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 23477 9367 23535 9373
rect 23477 9364 23489 9367
rect 23164 9336 23489 9364
rect 23164 9324 23170 9336
rect 23477 9333 23489 9336
rect 23523 9333 23535 9367
rect 29546 9364 29552 9376
rect 29507 9336 29552 9364
rect 23477 9327 23535 9333
rect 29546 9324 29552 9336
rect 29604 9324 29610 9376
rect 30190 9364 30196 9376
rect 30151 9336 30196 9364
rect 30190 9324 30196 9336
rect 30248 9324 30254 9376
rect 31110 9324 31116 9376
rect 31168 9364 31174 9376
rect 31573 9367 31631 9373
rect 31573 9364 31585 9367
rect 31168 9336 31585 9364
rect 31168 9324 31174 9336
rect 31573 9333 31585 9336
rect 31619 9333 31631 9367
rect 31573 9327 31631 9333
rect 32861 9367 32919 9373
rect 32861 9333 32873 9367
rect 32907 9364 32919 9367
rect 33428 9364 33456 9531
rect 33502 9528 33508 9580
rect 33560 9568 33566 9580
rect 33560 9540 33605 9568
rect 33560 9528 33566 9540
rect 33686 9528 33692 9580
rect 33744 9568 33750 9580
rect 34319 9569 34377 9575
rect 33744 9566 34284 9568
rect 34319 9566 34331 9569
rect 33744 9540 34331 9566
rect 33744 9528 33750 9540
rect 34256 9538 34331 9540
rect 34319 9535 34331 9538
rect 34365 9535 34377 9569
rect 34319 9529 34377 9535
rect 35526 9528 35532 9580
rect 35584 9568 35590 9580
rect 35713 9571 35771 9577
rect 35584 9540 35629 9568
rect 35584 9528 35590 9540
rect 35713 9537 35725 9571
rect 35759 9568 35771 9571
rect 36262 9568 36268 9580
rect 35759 9540 36268 9568
rect 35759 9537 35771 9540
rect 35713 9531 35771 9537
rect 36262 9528 36268 9540
rect 36320 9528 36326 9580
rect 37826 9528 37832 9580
rect 37884 9568 37890 9580
rect 37941 9571 37999 9577
rect 37941 9568 37953 9571
rect 37884 9540 37953 9568
rect 37884 9528 37890 9540
rect 37941 9537 37953 9540
rect 37987 9537 37999 9571
rect 37941 9531 37999 9537
rect 38120 9512 38148 9599
rect 41230 9596 41236 9608
rect 41288 9596 41294 9648
rect 45462 9636 45468 9648
rect 45423 9608 45468 9636
rect 45462 9596 45468 9608
rect 45520 9596 45526 9648
rect 45649 9639 45707 9645
rect 45649 9605 45661 9639
rect 45695 9636 45707 9639
rect 50249 9639 50307 9645
rect 50249 9636 50261 9639
rect 45695 9608 50261 9636
rect 45695 9605 45707 9608
rect 45649 9599 45707 9605
rect 50249 9605 50261 9608
rect 50295 9605 50307 9639
rect 53190 9636 53196 9648
rect 50249 9599 50307 9605
rect 52748 9608 53196 9636
rect 38189 9571 38247 9577
rect 38189 9537 38201 9571
rect 38235 9537 38247 9571
rect 38335 9571 38393 9577
rect 38335 9568 38347 9571
rect 38189 9531 38247 9537
rect 38328 9537 38347 9568
rect 38381 9537 38393 9571
rect 39117 9571 39175 9577
rect 39117 9568 39129 9571
rect 38328 9531 38393 9537
rect 38856 9540 39129 9568
rect 33778 9460 33784 9512
rect 33836 9500 33842 9512
rect 34149 9503 34207 9509
rect 34149 9500 34161 9503
rect 33836 9472 34161 9500
rect 33836 9460 33842 9472
rect 34149 9469 34161 9472
rect 34195 9500 34207 9503
rect 34195 9472 35572 9500
rect 34195 9469 34207 9472
rect 34149 9463 34207 9469
rect 35544 9444 35572 9472
rect 38102 9460 38108 9512
rect 38160 9460 38166 9512
rect 38212 9444 38240 9531
rect 38328 9500 38356 9531
rect 38856 9500 38884 9540
rect 39117 9537 39129 9540
rect 39163 9537 39175 9571
rect 40954 9568 40960 9580
rect 40915 9540 40960 9568
rect 39117 9531 39175 9537
rect 40954 9528 40960 9540
rect 41012 9528 41018 9580
rect 41138 9568 41144 9580
rect 41099 9540 41144 9568
rect 41138 9528 41144 9540
rect 41196 9528 41202 9580
rect 41322 9568 41328 9580
rect 41283 9540 41328 9568
rect 41322 9528 41328 9540
rect 41380 9528 41386 9580
rect 41506 9528 41512 9580
rect 41564 9568 41570 9580
rect 42613 9571 42671 9577
rect 42613 9568 42625 9571
rect 41564 9540 42625 9568
rect 41564 9528 41570 9540
rect 42613 9537 42625 9540
rect 42659 9537 42671 9571
rect 42613 9531 42671 9537
rect 45741 9571 45799 9577
rect 45741 9537 45753 9571
rect 45787 9537 45799 9571
rect 45741 9531 45799 9537
rect 38304 9472 38356 9500
rect 38488 9472 38884 9500
rect 33686 9432 33692 9444
rect 33647 9404 33692 9432
rect 33686 9392 33692 9404
rect 33744 9392 33750 9444
rect 35250 9432 35256 9444
rect 33796 9404 35256 9432
rect 33796 9364 33824 9404
rect 35250 9392 35256 9404
rect 35308 9392 35314 9444
rect 35526 9392 35532 9444
rect 35584 9392 35590 9444
rect 38194 9392 38200 9444
rect 38252 9392 38258 9444
rect 32907 9336 33824 9364
rect 32907 9333 32919 9336
rect 32861 9327 32919 9333
rect 34146 9324 34152 9376
rect 34204 9364 34210 9376
rect 34517 9367 34575 9373
rect 34517 9364 34529 9367
rect 34204 9336 34529 9364
rect 34204 9324 34210 9336
rect 34517 9333 34529 9336
rect 34563 9333 34575 9367
rect 34517 9327 34575 9333
rect 35342 9324 35348 9376
rect 35400 9364 35406 9376
rect 35897 9367 35955 9373
rect 35897 9364 35909 9367
rect 35400 9336 35909 9364
rect 35400 9324 35406 9336
rect 35897 9333 35909 9336
rect 35943 9364 35955 9367
rect 36170 9364 36176 9376
rect 35943 9336 36176 9364
rect 35943 9333 35955 9336
rect 35897 9327 35955 9333
rect 36170 9324 36176 9336
rect 36228 9324 36234 9376
rect 37550 9324 37556 9376
rect 37608 9364 37614 9376
rect 38304 9364 38332 9472
rect 38488 9441 38516 9472
rect 38930 9460 38936 9512
rect 38988 9500 38994 9512
rect 41966 9500 41972 9512
rect 38988 9472 41972 9500
rect 38988 9460 38994 9472
rect 41966 9460 41972 9472
rect 42024 9500 42030 9512
rect 42429 9503 42487 9509
rect 42429 9500 42441 9503
rect 42024 9472 42441 9500
rect 42024 9460 42030 9472
rect 42429 9469 42441 9472
rect 42475 9469 42487 9503
rect 45756 9500 45784 9531
rect 47026 9528 47032 9580
rect 47084 9568 47090 9580
rect 48222 9568 48228 9580
rect 47084 9540 48228 9568
rect 47084 9528 47090 9540
rect 48222 9528 48228 9540
rect 48280 9568 48286 9580
rect 48685 9571 48743 9577
rect 48685 9568 48697 9571
rect 48280 9540 48697 9568
rect 48280 9528 48286 9540
rect 48685 9537 48697 9540
rect 48731 9537 48743 9571
rect 48685 9531 48743 9537
rect 48869 9571 48927 9577
rect 48869 9537 48881 9571
rect 48915 9568 48927 9571
rect 49329 9571 49387 9577
rect 49329 9568 49341 9571
rect 48915 9540 49341 9568
rect 48915 9537 48927 9540
rect 48869 9531 48927 9537
rect 49329 9537 49341 9540
rect 49375 9568 49387 9571
rect 49970 9568 49976 9580
rect 49375 9540 49976 9568
rect 49375 9537 49387 9540
rect 49329 9531 49387 9537
rect 49970 9528 49976 9540
rect 50028 9528 50034 9580
rect 50893 9571 50951 9577
rect 50893 9537 50905 9571
rect 50939 9568 50951 9571
rect 51537 9571 51595 9577
rect 51537 9568 51549 9571
rect 50939 9540 51549 9568
rect 50939 9537 50951 9540
rect 50893 9531 50951 9537
rect 51537 9537 51549 9540
rect 51583 9568 51595 9571
rect 51810 9568 51816 9580
rect 51583 9540 51816 9568
rect 51583 9537 51595 9540
rect 51537 9531 51595 9537
rect 51810 9528 51816 9540
rect 51868 9528 51874 9580
rect 52748 9577 52776 9608
rect 53190 9596 53196 9608
rect 53248 9636 53254 9648
rect 53377 9639 53435 9645
rect 53377 9636 53389 9639
rect 53248 9608 53389 9636
rect 53248 9596 53254 9608
rect 53377 9605 53389 9608
rect 53423 9605 53435 9639
rect 56336 9636 56364 9667
rect 53377 9599 53435 9605
rect 53576 9608 56364 9636
rect 53576 9577 53604 9608
rect 52733 9571 52791 9577
rect 52733 9537 52745 9571
rect 52779 9537 52791 9571
rect 52733 9531 52791 9537
rect 52917 9571 52975 9577
rect 52917 9537 52929 9571
rect 52963 9568 52975 9571
rect 53561 9571 53619 9577
rect 53561 9568 53573 9571
rect 52963 9540 53573 9568
rect 52963 9537 52975 9540
rect 52917 9531 52975 9537
rect 53561 9537 53573 9540
rect 53607 9537 53619 9571
rect 53561 9531 53619 9537
rect 42429 9463 42487 9469
rect 43548 9472 45784 9500
rect 48501 9503 48559 9509
rect 38473 9435 38531 9441
rect 38473 9401 38485 9435
rect 38519 9401 38531 9435
rect 38473 9395 38531 9401
rect 39206 9392 39212 9444
rect 39264 9432 39270 9444
rect 43548 9432 43576 9472
rect 48501 9469 48513 9503
rect 48547 9500 48559 9503
rect 48590 9500 48596 9512
rect 48547 9472 48596 9500
rect 48547 9469 48559 9472
rect 48501 9463 48559 9469
rect 48590 9460 48596 9472
rect 48648 9460 48654 9512
rect 49510 9500 49516 9512
rect 49471 9472 49516 9500
rect 49510 9460 49516 9472
rect 49568 9460 49574 9512
rect 49602 9460 49608 9512
rect 49660 9500 49666 9512
rect 50433 9503 50491 9509
rect 50433 9500 50445 9503
rect 49660 9472 50445 9500
rect 49660 9460 49666 9472
rect 50433 9469 50445 9472
rect 50479 9469 50491 9503
rect 50433 9463 50491 9469
rect 50525 9503 50583 9509
rect 50525 9469 50537 9503
rect 50571 9469 50583 9503
rect 50525 9463 50583 9469
rect 50801 9503 50859 9509
rect 50801 9469 50813 9503
rect 50847 9469 50859 9503
rect 50801 9463 50859 9469
rect 39264 9404 43576 9432
rect 45465 9435 45523 9441
rect 39264 9392 39270 9404
rect 45465 9401 45477 9435
rect 45511 9432 45523 9435
rect 45554 9432 45560 9444
rect 45511 9404 45560 9432
rect 45511 9401 45523 9404
rect 45465 9395 45523 9401
rect 45554 9392 45560 9404
rect 45612 9392 45618 9444
rect 48608 9432 48636 9460
rect 50540 9432 50568 9463
rect 48608 9404 50568 9432
rect 50816 9432 50844 9463
rect 50982 9460 50988 9512
rect 51040 9500 51046 9512
rect 51353 9503 51411 9509
rect 51353 9500 51365 9503
rect 51040 9472 51365 9500
rect 51040 9460 51046 9472
rect 51353 9469 51365 9472
rect 51399 9469 51411 9503
rect 51353 9463 51411 9469
rect 51721 9503 51779 9509
rect 51721 9469 51733 9503
rect 51767 9500 51779 9503
rect 52748 9500 52776 9531
rect 51767 9472 52776 9500
rect 51767 9469 51779 9472
rect 51721 9463 51779 9469
rect 52932 9432 52960 9531
rect 54018 9528 54024 9580
rect 54076 9568 54082 9580
rect 54481 9571 54539 9577
rect 54481 9568 54493 9571
rect 54076 9540 54493 9568
rect 54076 9528 54082 9540
rect 54481 9537 54493 9540
rect 54527 9537 54539 9571
rect 55197 9571 55255 9577
rect 55197 9568 55209 9571
rect 54481 9531 54539 9537
rect 54864 9540 55209 9568
rect 50816 9404 52960 9432
rect 53558 9392 53564 9444
rect 53616 9432 53622 9444
rect 54297 9435 54355 9441
rect 53616 9404 54248 9432
rect 53616 9392 53622 9404
rect 41322 9364 41328 9376
rect 37608 9336 41328 9364
rect 37608 9324 37614 9336
rect 41322 9324 41328 9336
rect 41380 9324 41386 9376
rect 42797 9367 42855 9373
rect 42797 9333 42809 9367
rect 42843 9364 42855 9367
rect 45186 9364 45192 9376
rect 42843 9336 45192 9364
rect 42843 9333 42855 9336
rect 42797 9327 42855 9333
rect 45186 9324 45192 9336
rect 45244 9324 45250 9376
rect 52825 9367 52883 9373
rect 52825 9333 52837 9367
rect 52871 9364 52883 9367
rect 53006 9364 53012 9376
rect 52871 9336 53012 9364
rect 52871 9333 52883 9336
rect 52825 9327 52883 9333
rect 53006 9324 53012 9336
rect 53064 9324 53070 9376
rect 53742 9364 53748 9376
rect 53703 9336 53748 9364
rect 53742 9324 53748 9336
rect 53800 9324 53806 9376
rect 54220 9364 54248 9404
rect 54297 9401 54309 9435
rect 54343 9432 54355 9435
rect 54864 9432 54892 9540
rect 55197 9537 55209 9540
rect 55243 9537 55255 9571
rect 55197 9531 55255 9537
rect 54941 9503 54999 9509
rect 54941 9469 54953 9503
rect 54987 9469 54999 9503
rect 54941 9463 54999 9469
rect 54343 9404 54892 9432
rect 54343 9401 54355 9404
rect 54297 9395 54355 9401
rect 54956 9364 54984 9463
rect 54220 9336 54984 9364
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 9490 9160 9496 9172
rect 4264 9132 9496 9160
rect 4264 9092 4292 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 10962 9160 10968 9172
rect 9600 9132 10548 9160
rect 10923 9132 10968 9160
rect 1688 9064 4292 9092
rect 1688 9033 1716 9064
rect 4338 9052 4344 9104
rect 4396 9092 4402 9104
rect 9600 9092 9628 9132
rect 4396 9064 9628 9092
rect 10520 9092 10548 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 11756 9132 17601 9160
rect 11756 9120 11762 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 20070 9160 20076 9172
rect 17920 9132 18092 9160
rect 20031 9132 20076 9160
rect 17920 9120 17926 9132
rect 16666 9092 16672 9104
rect 10520 9064 16672 9092
rect 4396 9052 4402 9064
rect 16666 9052 16672 9064
rect 16724 9052 16730 9104
rect 17310 9092 17316 9104
rect 17052 9064 17316 9092
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 9490 9024 9496 9036
rect 1673 8987 1731 8993
rect 7208 8996 9496 9024
rect 1394 8956 1400 8968
rect 1355 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 4246 8956 4252 8968
rect 4207 8928 4252 8956
rect 3973 8919 4031 8925
rect 3988 8888 4016 8919
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 7208 8965 7236 8996
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 14277 9027 14335 9033
rect 14277 9024 14289 9027
rect 13964 8996 14289 9024
rect 13964 8984 13970 8996
rect 14277 8993 14289 8996
rect 14323 9024 14335 9027
rect 14642 9024 14648 9036
rect 14323 8996 14648 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 17052 9033 17080 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 17604 9064 18000 9092
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16632 8996 16957 9024
rect 16632 8984 16638 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 16945 8987 17003 8993
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 17126 8984 17132 9036
rect 17184 9024 17190 9036
rect 17604 9024 17632 9064
rect 17770 9024 17776 9036
rect 17184 8996 17632 9024
rect 17731 8996 17776 9024
rect 17184 8984 17190 8996
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 17972 9033 18000 9064
rect 18064 9033 18092 9132
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 22428 9132 22569 9160
rect 22428 9120 22434 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 25869 9163 25927 9169
rect 25869 9129 25881 9163
rect 25915 9160 25927 9163
rect 26326 9160 26332 9172
rect 25915 9132 26332 9160
rect 25915 9129 25927 9132
rect 25869 9123 25927 9129
rect 26326 9120 26332 9132
rect 26384 9120 26390 9172
rect 31849 9163 31907 9169
rect 26436 9132 31754 9160
rect 21358 9092 21364 9104
rect 20272 9064 21364 9092
rect 20272 9033 20300 9064
rect 21358 9052 21364 9064
rect 21416 9092 21422 9104
rect 21416 9064 22094 9092
rect 21416 9052 21422 9064
rect 17957 9027 18015 9033
rect 17957 8993 17969 9027
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 20257 9027 20315 9033
rect 20257 8993 20269 9027
rect 20303 8993 20315 9027
rect 20622 9024 20628 9036
rect 20583 8996 20628 9024
rect 20257 8987 20315 8993
rect 20622 8984 20628 8996
rect 20680 8984 20686 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20732 8996 21281 9024
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 7193 8919 7251 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 9582 8956 9588 8968
rect 9543 8928 9588 8956
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9841 8959 9899 8965
rect 9841 8956 9853 8959
rect 9732 8928 9853 8956
rect 9732 8916 9738 8928
rect 9841 8925 9853 8928
rect 9887 8925 9899 8959
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 9841 8919 9899 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 14366 8956 14372 8968
rect 12575 8928 14372 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 11698 8888 11704 8900
rect 3988 8860 11704 8888
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 3786 8820 3792 8832
rect 3747 8792 3792 8820
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 4120 8792 4169 8820
rect 4120 8780 4126 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 7006 8820 7012 8832
rect 6967 8792 7012 8820
rect 4157 8783 4215 8789
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 12544 8820 12572 8919
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14476 8888 14504 8919
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 16758 8956 16764 8968
rect 14608 8928 14653 8956
rect 16719 8928 16764 8956
rect 14608 8916 14614 8928
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 16850 8916 16856 8968
rect 16908 8956 16914 8968
rect 17218 8956 17224 8968
rect 16908 8928 17224 8956
rect 16908 8927 16988 8928
rect 16908 8916 16914 8927
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 20349 8959 20407 8965
rect 17920 8928 17965 8956
rect 17920 8916 17926 8928
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20732 8956 20760 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 22066 9024 22094 9064
rect 23566 9052 23572 9104
rect 23624 9092 23630 9104
rect 26436 9092 26464 9132
rect 23624 9064 26464 9092
rect 23624 9052 23630 9064
rect 22741 9027 22799 9033
rect 22741 9024 22753 9027
rect 22066 8996 22753 9024
rect 21269 8987 21327 8993
rect 22741 8993 22753 8996
rect 22787 8993 22799 9027
rect 23750 9024 23756 9036
rect 22741 8987 22799 8993
rect 22848 8996 23756 9024
rect 20395 8928 20760 8956
rect 21177 8959 21235 8965
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 20640 8900 20668 8928
rect 21177 8925 21189 8959
rect 21223 8925 21235 8959
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21177 8919 21235 8925
rect 14476 8860 18276 8888
rect 10560 8792 12572 8820
rect 14093 8823 14151 8829
rect 10560 8780 10566 8792
rect 14093 8789 14105 8823
rect 14139 8820 14151 8823
rect 14182 8820 14188 8832
rect 14139 8792 14188 8820
rect 14139 8789 14151 8792
rect 14093 8783 14151 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 16577 8823 16635 8829
rect 16577 8820 16589 8823
rect 15804 8792 16589 8820
rect 15804 8780 15810 8792
rect 16577 8789 16589 8792
rect 16623 8789 16635 8823
rect 18248 8820 18276 8860
rect 20622 8848 20628 8900
rect 20680 8848 20686 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 21192 8888 21220 8919
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 22848 8965 22876 8996
rect 23750 8984 23756 8996
rect 23808 8984 23814 9036
rect 25593 9027 25651 9033
rect 25593 8993 25605 9027
rect 25639 9024 25651 9027
rect 26050 9024 26056 9036
rect 25639 8996 26056 9024
rect 25639 8993 25651 8996
rect 25593 8987 25651 8993
rect 26050 8984 26056 8996
rect 26108 8984 26114 9036
rect 26878 8984 26884 9036
rect 26936 9024 26942 9036
rect 31726 9024 31754 9132
rect 31849 9129 31861 9163
rect 31895 9160 31907 9163
rect 32306 9160 32312 9172
rect 31895 9132 32312 9160
rect 31895 9129 31907 9132
rect 31849 9123 31907 9129
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 33502 9120 33508 9172
rect 33560 9160 33566 9172
rect 35437 9163 35495 9169
rect 35437 9160 35449 9163
rect 33560 9132 35449 9160
rect 33560 9120 33566 9132
rect 35437 9129 35449 9132
rect 35483 9160 35495 9163
rect 37550 9160 37556 9172
rect 35483 9132 37556 9160
rect 35483 9129 35495 9132
rect 35437 9123 35495 9129
rect 37550 9120 37556 9132
rect 37608 9120 37614 9172
rect 40034 9160 40040 9172
rect 37660 9132 40040 9160
rect 34330 9052 34336 9104
rect 34388 9092 34394 9104
rect 36357 9095 36415 9101
rect 36357 9092 36369 9095
rect 34388 9064 36369 9092
rect 34388 9052 34394 9064
rect 36357 9061 36369 9064
rect 36403 9092 36415 9095
rect 37660 9092 37688 9132
rect 40034 9120 40040 9132
rect 40092 9120 40098 9172
rect 41414 9120 41420 9172
rect 41472 9160 41478 9172
rect 41785 9163 41843 9169
rect 41785 9160 41797 9163
rect 41472 9132 41797 9160
rect 41472 9120 41478 9132
rect 41785 9129 41797 9132
rect 41831 9129 41843 9163
rect 41785 9123 41843 9129
rect 50706 9120 50712 9172
rect 50764 9160 50770 9172
rect 52273 9163 52331 9169
rect 52273 9160 52285 9163
rect 50764 9132 52285 9160
rect 50764 9120 50770 9132
rect 52273 9129 52285 9132
rect 52319 9129 52331 9163
rect 52273 9123 52331 9129
rect 53006 9120 53012 9172
rect 53064 9160 53070 9172
rect 53837 9163 53895 9169
rect 53837 9160 53849 9163
rect 53064 9132 53849 9160
rect 53064 9120 53070 9132
rect 53837 9129 53849 9132
rect 53883 9129 53895 9163
rect 54018 9160 54024 9172
rect 53979 9132 54024 9160
rect 53837 9123 53895 9129
rect 54018 9120 54024 9132
rect 54076 9120 54082 9172
rect 36403 9064 37688 9092
rect 36403 9061 36415 9064
rect 36357 9055 36415 9061
rect 39114 9052 39120 9104
rect 39172 9092 39178 9104
rect 39172 9064 41414 9092
rect 39172 9052 39178 9064
rect 32398 9024 32404 9036
rect 26936 8996 30144 9024
rect 31726 8996 32404 9024
rect 26936 8984 26942 8996
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 23661 8959 23719 8965
rect 23661 8956 23673 8959
rect 22833 8919 22891 8925
rect 22940 8928 23673 8956
rect 21726 8888 21732 8900
rect 20772 8860 20817 8888
rect 21192 8860 21732 8888
rect 20772 8848 20778 8860
rect 21726 8848 21732 8860
rect 21784 8888 21790 8900
rect 22940 8888 22968 8928
rect 23661 8925 23673 8928
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24578 8956 24584 8968
rect 23891 8928 24584 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 25501 8959 25559 8965
rect 25501 8925 25513 8959
rect 25547 8956 25559 8959
rect 26234 8956 26240 8968
rect 25547 8928 26240 8956
rect 25547 8925 25559 8928
rect 25501 8919 25559 8925
rect 26234 8916 26240 8928
rect 26292 8916 26298 8968
rect 28166 8916 28172 8968
rect 28224 8956 28230 8968
rect 30006 8956 30012 8968
rect 28224 8928 30012 8956
rect 28224 8916 28230 8928
rect 30006 8916 30012 8928
rect 30064 8916 30070 8968
rect 30116 8956 30144 8996
rect 32398 8984 32404 8996
rect 32456 8984 32462 9036
rect 32493 9027 32551 9033
rect 32493 8993 32505 9027
rect 32539 9024 32551 9027
rect 33686 9024 33692 9036
rect 32539 8996 33692 9024
rect 32539 8993 32551 8996
rect 32493 8987 32551 8993
rect 33686 8984 33692 8996
rect 33744 8984 33750 9036
rect 35894 8984 35900 9036
rect 35952 9024 35958 9036
rect 36814 9024 36820 9036
rect 35952 8996 36820 9024
rect 35952 8984 35958 8996
rect 36814 8984 36820 8996
rect 36872 8984 36878 9036
rect 41386 9024 41414 9064
rect 42150 9052 42156 9104
rect 42208 9092 42214 9104
rect 46934 9092 46940 9104
rect 42208 9064 46940 9092
rect 42208 9052 42214 9064
rect 46934 9052 46940 9064
rect 46992 9052 46998 9104
rect 50154 9092 50160 9104
rect 50115 9064 50160 9092
rect 50154 9052 50160 9064
rect 50212 9052 50218 9104
rect 42429 9027 42487 9033
rect 42429 9024 42441 9027
rect 41386 8996 42441 9024
rect 42429 8993 42441 8996
rect 42475 9024 42487 9027
rect 42518 9024 42524 9036
rect 42475 8996 42524 9024
rect 42475 8993 42487 8996
rect 42429 8987 42487 8993
rect 42518 8984 42524 8996
rect 42576 8984 42582 9036
rect 47026 9024 47032 9036
rect 45020 8996 47032 9024
rect 30116 8928 34100 8956
rect 23106 8888 23112 8900
rect 21784 8860 22968 8888
rect 23067 8860 23112 8888
rect 21784 8848 21790 8860
rect 23106 8848 23112 8860
rect 23164 8848 23170 8900
rect 23198 8848 23204 8900
rect 23256 8888 23262 8900
rect 30276 8891 30334 8897
rect 23256 8860 23301 8888
rect 23256 8848 23262 8860
rect 30276 8857 30288 8891
rect 30322 8888 30334 8891
rect 30926 8888 30932 8900
rect 30322 8860 30932 8888
rect 30322 8857 30334 8860
rect 30276 8851 30334 8857
rect 30926 8848 30932 8860
rect 30984 8848 30990 8900
rect 32217 8891 32275 8897
rect 32217 8888 32229 8891
rect 31726 8860 32229 8888
rect 23124 8820 23152 8848
rect 18248 8792 23152 8820
rect 16577 8783 16635 8789
rect 30834 8780 30840 8832
rect 30892 8820 30898 8832
rect 31389 8823 31447 8829
rect 31389 8820 31401 8823
rect 30892 8792 31401 8820
rect 30892 8780 30898 8792
rect 31389 8789 31401 8792
rect 31435 8820 31447 8823
rect 31726 8820 31754 8860
rect 32217 8857 32229 8860
rect 32263 8857 32275 8891
rect 32217 8851 32275 8857
rect 32490 8848 32496 8900
rect 32548 8888 32554 8900
rect 33594 8888 33600 8900
rect 32548 8860 33600 8888
rect 32548 8848 32554 8860
rect 33594 8848 33600 8860
rect 33652 8848 33658 8900
rect 31435 8792 31754 8820
rect 31435 8789 31447 8792
rect 31389 8783 31447 8789
rect 32030 8780 32036 8832
rect 32088 8820 32094 8832
rect 32309 8823 32367 8829
rect 32309 8820 32321 8823
rect 32088 8792 32321 8820
rect 32088 8780 32094 8792
rect 32309 8789 32321 8792
rect 32355 8789 32367 8823
rect 33962 8820 33968 8832
rect 33923 8792 33968 8820
rect 32309 8783 32367 8789
rect 33962 8780 33968 8792
rect 34020 8780 34026 8832
rect 34072 8820 34100 8928
rect 34146 8916 34152 8968
rect 34204 8956 34210 8968
rect 35342 8956 35348 8968
rect 34204 8928 34249 8956
rect 35303 8928 35348 8956
rect 34204 8916 34210 8928
rect 35342 8916 35348 8928
rect 35400 8916 35406 8968
rect 37918 8956 37924 8968
rect 35452 8928 36216 8956
rect 37879 8928 37924 8956
rect 34330 8848 34336 8900
rect 34388 8888 34394 8900
rect 35452 8888 35480 8928
rect 34388 8860 35480 8888
rect 36081 8891 36139 8897
rect 34388 8848 34394 8860
rect 36081 8857 36093 8891
rect 36127 8857 36139 8891
rect 36188 8888 36216 8928
rect 37918 8916 37924 8928
rect 37976 8916 37982 8968
rect 38010 8916 38016 8968
rect 38068 8956 38074 8968
rect 38177 8959 38235 8965
rect 38177 8956 38189 8959
rect 38068 8928 38189 8956
rect 38068 8916 38074 8928
rect 38177 8925 38189 8928
rect 38223 8925 38235 8959
rect 45020 8956 45048 8996
rect 47026 8984 47032 8996
rect 47084 8984 47090 9036
rect 45186 8956 45192 8968
rect 38177 8919 38235 8925
rect 38304 8928 45048 8956
rect 45147 8928 45192 8956
rect 38304 8888 38332 8928
rect 45186 8916 45192 8928
rect 45244 8916 45250 8968
rect 50062 8916 50068 8968
rect 50120 8956 50126 8968
rect 50341 8959 50399 8965
rect 50341 8956 50353 8959
rect 50120 8928 50353 8956
rect 50120 8916 50126 8928
rect 50341 8925 50353 8928
rect 50387 8925 50399 8959
rect 50341 8919 50399 8925
rect 50433 8959 50491 8965
rect 50433 8925 50445 8959
rect 50479 8956 50491 8959
rect 50706 8956 50712 8968
rect 50479 8928 50712 8956
rect 50479 8925 50491 8928
rect 50433 8919 50491 8925
rect 50706 8916 50712 8928
rect 50764 8956 50770 8968
rect 50982 8956 50988 8968
rect 50764 8928 50988 8956
rect 50764 8916 50770 8928
rect 50982 8916 50988 8928
rect 51040 8916 51046 8968
rect 52181 8959 52239 8965
rect 52181 8925 52193 8959
rect 52227 8956 52239 8959
rect 53282 8956 53288 8968
rect 52227 8928 53288 8956
rect 52227 8925 52239 8928
rect 52181 8919 52239 8925
rect 53282 8916 53288 8928
rect 53340 8916 53346 8968
rect 50157 8891 50215 8897
rect 50157 8888 50169 8891
rect 36188 8860 38332 8888
rect 38396 8860 50169 8888
rect 36081 8851 36139 8857
rect 34698 8820 34704 8832
rect 34072 8792 34704 8820
rect 34698 8780 34704 8792
rect 34756 8820 34762 8832
rect 36096 8820 36124 8851
rect 34756 8792 36124 8820
rect 34756 8780 34762 8792
rect 36538 8780 36544 8832
rect 36596 8820 36602 8832
rect 38396 8820 38424 8860
rect 50157 8857 50169 8860
rect 50203 8888 50215 8891
rect 53650 8888 53656 8900
rect 50203 8860 51074 8888
rect 53611 8860 53656 8888
rect 50203 8857 50215 8860
rect 50157 8851 50215 8857
rect 39298 8820 39304 8832
rect 36596 8792 38424 8820
rect 39259 8792 39304 8820
rect 36596 8780 36602 8792
rect 39298 8780 39304 8792
rect 39356 8780 39362 8832
rect 39390 8780 39396 8832
rect 39448 8820 39454 8832
rect 42150 8820 42156 8832
rect 39448 8792 42156 8820
rect 39448 8780 39454 8792
rect 42150 8780 42156 8792
rect 42208 8780 42214 8832
rect 42245 8823 42303 8829
rect 42245 8789 42257 8823
rect 42291 8820 42303 8823
rect 42610 8820 42616 8832
rect 42291 8792 42616 8820
rect 42291 8789 42303 8792
rect 42245 8783 42303 8789
rect 42610 8780 42616 8792
rect 42668 8780 42674 8832
rect 45002 8820 45008 8832
rect 44963 8792 45008 8820
rect 45002 8780 45008 8792
rect 45060 8780 45066 8832
rect 51046 8820 51074 8860
rect 53650 8848 53656 8860
rect 53708 8848 53714 8900
rect 53742 8848 53748 8900
rect 53800 8888 53806 8900
rect 53853 8891 53911 8897
rect 53853 8888 53865 8891
rect 53800 8860 53865 8888
rect 53800 8848 53806 8860
rect 53853 8857 53865 8860
rect 53899 8857 53911 8891
rect 53853 8851 53911 8857
rect 52914 8820 52920 8832
rect 51046 8792 52920 8820
rect 52914 8780 52920 8792
rect 52972 8780 52978 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 2041 8619 2099 8625
rect 2041 8585 2053 8619
rect 2087 8616 2099 8619
rect 4338 8616 4344 8628
rect 2087 8588 4344 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 7374 8616 7380 8628
rect 4448 8588 7380 8616
rect 1762 8548 1768 8560
rect 1723 8520 1768 8548
rect 1762 8508 1768 8520
rect 1820 8508 1826 8560
rect 2860 8551 2918 8557
rect 2860 8517 2872 8551
rect 2906 8548 2918 8551
rect 3786 8548 3792 8560
rect 2906 8520 3792 8548
rect 2906 8517 2918 8520
rect 2860 8511 2918 8517
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 4448 8548 4476 8588
rect 7374 8576 7380 8588
rect 7432 8616 7438 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7432 8588 7757 8616
rect 7432 8576 7438 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9858 8616 9864 8628
rect 9723 8588 9864 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10502 8616 10508 8628
rect 10091 8588 10508 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 11756 8588 16681 8616
rect 11756 8576 11762 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 16908 8588 17264 8616
rect 16908 8576 16914 8588
rect 4028 8520 4476 8548
rect 6632 8551 6690 8557
rect 4028 8508 4034 8520
rect 6632 8517 6644 8551
rect 6678 8548 6690 8551
rect 7006 8548 7012 8560
rect 6678 8520 7012 8548
rect 6678 8517 6690 8520
rect 6632 8511 6690 8517
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 13446 8548 13452 8560
rect 7576 8520 13452 8548
rect 2222 8440 2228 8492
rect 2280 8480 2286 8492
rect 2280 8452 4200 8480
rect 2280 8440 2286 8452
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2096 8384 2605 8412
rect 2096 8372 2102 8384
rect 2593 8381 2605 8384
rect 2639 8381 2651 8415
rect 2593 8375 2651 8381
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4062 8344 4068 8356
rect 4019 8316 4068 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4172 8344 4200 8452
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 4614 8480 4620 8492
rect 4304 8452 4620 8480
rect 4304 8440 4310 8452
rect 4614 8440 4620 8452
rect 4672 8480 4678 8492
rect 7466 8480 7472 8492
rect 4672 8452 7472 8480
rect 4672 8440 4678 8452
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 6362 8412 6368 8424
rect 6323 8384 6368 8412
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 7576 8344 7604 8520
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 14550 8508 14556 8560
rect 14608 8548 14614 8560
rect 14608 8520 15608 8548
rect 14608 8508 14614 8520
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9548 8452 11468 8480
rect 9548 8440 9554 8452
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 8352 8384 10149 8412
rect 8352 8372 8358 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10137 8375 10195 8381
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10686 8412 10692 8424
rect 10367 8384 10692 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 11440 8412 11468 8452
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 12768 8452 13185 8480
rect 12768 8440 12774 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13354 8480 13360 8492
rect 13311 8452 13360 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8480 13783 8483
rect 13814 8480 13820 8492
rect 13771 8452 13820 8480
rect 13771 8449 13783 8452
rect 13725 8443 13783 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14461 8483 14519 8489
rect 14240 8452 14412 8480
rect 14240 8440 14246 8452
rect 14384 8421 14412 8452
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14734 8480 14740 8492
rect 14507 8452 14740 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 14369 8415 14427 8421
rect 11440 8384 14320 8412
rect 12986 8344 12992 8356
rect 4172 8316 6408 8344
rect 6380 8276 6408 8316
rect 7300 8316 7604 8344
rect 12947 8316 12992 8344
rect 7300 8276 7328 8316
rect 12986 8304 12992 8316
rect 13044 8304 13050 8356
rect 13078 8304 13084 8356
rect 13136 8344 13142 8356
rect 14185 8347 14243 8353
rect 14185 8344 14197 8347
rect 13136 8316 14197 8344
rect 13136 8304 13142 8316
rect 14185 8313 14197 8316
rect 14231 8313 14243 8347
rect 14292 8344 14320 8384
rect 14369 8381 14381 8415
rect 14415 8381 14427 8415
rect 14550 8412 14556 8424
rect 14511 8384 14556 8412
rect 14369 8375 14427 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 15470 8412 15476 8424
rect 14691 8384 15476 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15580 8412 15608 8520
rect 15654 8508 15660 8560
rect 15712 8548 15718 8560
rect 16758 8548 16764 8560
rect 15712 8520 16764 8548
rect 15712 8508 15718 8520
rect 16758 8508 16764 8520
rect 16816 8548 16822 8560
rect 17126 8548 17132 8560
rect 16816 8520 17132 8548
rect 16816 8508 16822 8520
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17236 8548 17264 8588
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 22094 8616 22100 8628
rect 20772 8588 22100 8616
rect 20772 8576 20778 8588
rect 22094 8576 22100 8588
rect 22152 8616 22158 8628
rect 23198 8616 23204 8628
rect 22152 8588 23204 8616
rect 22152 8576 22158 8588
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 30926 8616 30932 8628
rect 30887 8588 30932 8616
rect 30926 8576 30932 8588
rect 30984 8576 30990 8628
rect 31018 8576 31024 8628
rect 31076 8616 31082 8628
rect 31076 8588 31754 8616
rect 31076 8576 31082 8588
rect 24578 8548 24584 8560
rect 17236 8520 24584 8548
rect 24578 8508 24584 8520
rect 24636 8508 24642 8560
rect 27798 8508 27804 8560
rect 27856 8548 27862 8560
rect 28077 8551 28135 8557
rect 28077 8548 28089 8551
rect 27856 8520 28089 8548
rect 27856 8508 27862 8520
rect 28077 8517 28089 8520
rect 28123 8517 28135 8551
rect 28077 8511 28135 8517
rect 28166 8508 28172 8560
rect 28224 8548 28230 8560
rect 28293 8551 28351 8557
rect 28293 8548 28305 8551
rect 28224 8520 28305 8548
rect 28224 8508 28230 8520
rect 28293 8517 28305 8520
rect 28339 8548 28351 8551
rect 31726 8548 31754 8588
rect 34330 8576 34336 8628
rect 34388 8616 34394 8628
rect 36538 8616 36544 8628
rect 34388 8588 36544 8616
rect 34388 8576 34394 8588
rect 36538 8576 36544 8588
rect 36596 8576 36602 8628
rect 38102 8576 38108 8628
rect 38160 8616 38166 8628
rect 38565 8619 38623 8625
rect 38565 8616 38577 8619
rect 38160 8588 38577 8616
rect 38160 8576 38166 8588
rect 38565 8585 38577 8588
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 39025 8619 39083 8625
rect 39025 8585 39037 8619
rect 39071 8616 39083 8619
rect 39390 8616 39396 8628
rect 39071 8588 39396 8616
rect 39071 8585 39083 8588
rect 39025 8579 39083 8585
rect 39390 8576 39396 8588
rect 39448 8576 39454 8628
rect 40862 8616 40868 8628
rect 39500 8588 40868 8616
rect 28339 8520 31248 8548
rect 31726 8520 33916 8548
rect 28339 8517 28351 8520
rect 28293 8511 28351 8517
rect 15746 8480 15752 8492
rect 15707 8452 15752 8480
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16206 8480 16212 8492
rect 15887 8452 16212 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16942 8440 16948 8492
rect 17000 8480 17006 8492
rect 23566 8480 23572 8492
rect 17000 8452 17045 8480
rect 23527 8452 23572 8480
rect 17000 8440 17006 8452
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 23750 8480 23756 8492
rect 23707 8452 23756 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15580 8384 15945 8412
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16025 8415 16083 8421
rect 16025 8381 16037 8415
rect 16071 8412 16083 8415
rect 16666 8412 16672 8424
rect 16071 8384 16672 8412
rect 16071 8381 16083 8384
rect 16025 8375 16083 8381
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 14292 8316 15577 8344
rect 14185 8307 14243 8313
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 15948 8344 15976 8375
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 16850 8412 16856 8424
rect 16811 8384 16856 8412
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17034 8412 17040 8424
rect 16947 8384 17040 8412
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 17126 8372 17132 8424
rect 17184 8412 17190 8424
rect 17586 8412 17592 8424
rect 17184 8384 17592 8412
rect 17184 8372 17190 8384
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 23842 8412 23848 8424
rect 23803 8384 23848 8412
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 27448 8412 27476 8443
rect 27522 8440 27528 8492
rect 27580 8480 27586 8492
rect 27617 8483 27675 8489
rect 27617 8480 27629 8483
rect 27580 8452 27629 8480
rect 27580 8440 27586 8452
rect 27617 8449 27629 8452
rect 27663 8480 27675 8483
rect 31110 8480 31116 8492
rect 27663 8452 28488 8480
rect 31071 8452 31116 8480
rect 27663 8449 27675 8452
rect 27617 8443 27675 8449
rect 28074 8412 28080 8424
rect 27448 8384 28080 8412
rect 28074 8372 28080 8384
rect 28132 8372 28138 8424
rect 17052 8344 17080 8372
rect 21358 8344 21364 8356
rect 15948 8316 17080 8344
rect 19306 8316 21364 8344
rect 15565 8307 15623 8313
rect 6380 8248 7328 8276
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 19306 8276 19334 8316
rect 21358 8304 21364 8316
rect 21416 8344 21422 8356
rect 21726 8344 21732 8356
rect 21416 8316 21732 8344
rect 21416 8304 21422 8316
rect 21726 8304 21732 8316
rect 21784 8304 21790 8356
rect 28460 8353 28488 8452
rect 31110 8440 31116 8452
rect 31168 8440 31174 8492
rect 31220 8480 31248 8520
rect 33778 8480 33784 8492
rect 31220 8452 33784 8480
rect 33778 8440 33784 8452
rect 33836 8440 33842 8492
rect 33888 8480 33916 8520
rect 33962 8508 33968 8560
rect 34020 8548 34026 8560
rect 34118 8551 34176 8557
rect 34118 8548 34130 8551
rect 34020 8520 34130 8548
rect 34020 8508 34026 8520
rect 34118 8517 34130 8520
rect 34164 8517 34176 8551
rect 34118 8511 34176 8517
rect 35802 8508 35808 8560
rect 35860 8548 35866 8560
rect 39500 8548 39528 8588
rect 40862 8576 40868 8588
rect 40920 8576 40926 8628
rect 41138 8576 41144 8628
rect 41196 8616 41202 8628
rect 42429 8619 42487 8625
rect 42429 8616 42441 8619
rect 41196 8588 42441 8616
rect 41196 8576 41202 8588
rect 42429 8585 42441 8588
rect 42475 8585 42487 8619
rect 42429 8579 42487 8585
rect 50062 8576 50068 8628
rect 50120 8616 50126 8628
rect 50614 8616 50620 8628
rect 50120 8588 50620 8616
rect 50120 8576 50126 8588
rect 50614 8576 50620 8588
rect 50672 8616 50678 8628
rect 50709 8619 50767 8625
rect 50709 8616 50721 8619
rect 50672 8588 50721 8616
rect 50672 8576 50678 8588
rect 50709 8585 50721 8588
rect 50755 8585 50767 8619
rect 50709 8579 50767 8585
rect 35860 8520 39528 8548
rect 35860 8508 35866 8520
rect 40034 8508 40040 8560
rect 40092 8548 40098 8560
rect 40313 8551 40371 8557
rect 40313 8548 40325 8551
rect 40092 8520 40325 8548
rect 40092 8508 40098 8520
rect 40313 8517 40325 8520
rect 40359 8548 40371 8551
rect 40770 8548 40776 8560
rect 40359 8520 40776 8548
rect 40359 8517 40371 8520
rect 40313 8511 40371 8517
rect 40770 8508 40776 8520
rect 40828 8508 40834 8560
rect 42518 8508 42524 8560
rect 42576 8548 42582 8560
rect 42576 8520 43024 8548
rect 42576 8508 42582 8520
rect 36081 8483 36139 8489
rect 33888 8452 35664 8480
rect 30006 8372 30012 8424
rect 30064 8412 30070 8424
rect 33873 8415 33931 8421
rect 33873 8412 33885 8415
rect 30064 8384 33885 8412
rect 30064 8372 30070 8384
rect 33873 8381 33885 8384
rect 33919 8381 33931 8415
rect 33873 8375 33931 8381
rect 28445 8347 28503 8353
rect 28445 8313 28457 8347
rect 28491 8313 28503 8347
rect 28445 8307 28503 8313
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 35636 8344 35664 8452
rect 36081 8449 36093 8483
rect 36127 8480 36139 8483
rect 36170 8480 36176 8492
rect 36127 8452 36176 8480
rect 36127 8449 36139 8452
rect 36081 8443 36139 8449
rect 36170 8440 36176 8452
rect 36228 8440 36234 8492
rect 36262 8440 36268 8492
rect 36320 8480 36326 8492
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 36320 8452 37473 8480
rect 36320 8440 36326 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8480 38991 8483
rect 39298 8480 39304 8492
rect 38979 8452 39304 8480
rect 38979 8449 38991 8452
rect 38933 8443 38991 8449
rect 35802 8372 35808 8424
rect 35860 8412 35866 8424
rect 38948 8412 38976 8443
rect 39298 8440 39304 8452
rect 39356 8440 39362 8492
rect 40126 8480 40132 8492
rect 40087 8452 40132 8480
rect 40126 8440 40132 8452
rect 40184 8440 40190 8492
rect 40218 8440 40224 8492
rect 40276 8480 40282 8492
rect 40494 8489 40500 8492
rect 40451 8483 40500 8489
rect 40276 8452 40321 8480
rect 40276 8440 40282 8452
rect 40451 8449 40463 8483
rect 40497 8449 40500 8483
rect 40451 8443 40500 8449
rect 40494 8440 40500 8443
rect 40552 8440 40558 8492
rect 42794 8480 42800 8492
rect 42755 8452 42800 8480
rect 42794 8440 42800 8452
rect 42852 8440 42858 8492
rect 39114 8412 39120 8424
rect 35860 8384 38976 8412
rect 39075 8384 39120 8412
rect 35860 8372 35866 8384
rect 39114 8372 39120 8384
rect 39172 8372 39178 8424
rect 40589 8415 40647 8421
rect 40589 8412 40601 8415
rect 39224 8384 40601 8412
rect 39224 8344 39252 8384
rect 40589 8381 40601 8384
rect 40635 8381 40647 8415
rect 42242 8412 42248 8424
rect 40589 8375 40647 8381
rect 40788 8384 42248 8412
rect 30340 8316 33916 8344
rect 35636 8316 39252 8344
rect 39945 8347 40003 8353
rect 30340 8304 30346 8316
rect 13504 8248 19334 8276
rect 13504 8236 13510 8248
rect 23750 8236 23756 8288
rect 23808 8276 23814 8288
rect 23808 8248 23853 8276
rect 23808 8236 23814 8248
rect 27154 8236 27160 8288
rect 27212 8276 27218 8288
rect 27433 8279 27491 8285
rect 27433 8276 27445 8279
rect 27212 8248 27445 8276
rect 27212 8236 27218 8248
rect 27433 8245 27445 8248
rect 27479 8245 27491 8279
rect 27433 8239 27491 8245
rect 28261 8279 28319 8285
rect 28261 8245 28273 8279
rect 28307 8276 28319 8279
rect 30190 8276 30196 8288
rect 28307 8248 30196 8276
rect 28307 8245 28319 8248
rect 28261 8239 28319 8245
rect 30190 8236 30196 8248
rect 30248 8236 30254 8288
rect 31386 8236 31392 8288
rect 31444 8276 31450 8288
rect 33410 8276 33416 8288
rect 31444 8248 33416 8276
rect 31444 8236 31450 8248
rect 33410 8236 33416 8248
rect 33468 8236 33474 8288
rect 33888 8276 33916 8316
rect 39945 8313 39957 8347
rect 39991 8344 40003 8347
rect 40034 8344 40040 8356
rect 39991 8316 40040 8344
rect 39991 8313 40003 8316
rect 39945 8307 40003 8313
rect 40034 8304 40040 8316
rect 40092 8304 40098 8356
rect 40126 8304 40132 8356
rect 40184 8344 40190 8356
rect 40788 8344 40816 8384
rect 42242 8372 42248 8384
rect 42300 8372 42306 8424
rect 42996 8421 43024 8520
rect 45002 8508 45008 8560
rect 45060 8548 45066 8560
rect 45710 8551 45768 8557
rect 45710 8548 45722 8551
rect 45060 8520 45722 8548
rect 45060 8508 45066 8520
rect 45710 8517 45722 8520
rect 45756 8517 45768 8551
rect 52638 8548 52644 8560
rect 45710 8511 45768 8517
rect 49344 8520 52644 8548
rect 43714 8440 43720 8492
rect 43772 8480 43778 8492
rect 45465 8483 45523 8489
rect 45465 8480 45477 8483
rect 43772 8452 45477 8480
rect 43772 8440 43778 8452
rect 45465 8449 45477 8452
rect 45511 8480 45523 8483
rect 45554 8480 45560 8492
rect 45511 8452 45560 8480
rect 45511 8449 45523 8452
rect 45465 8443 45523 8449
rect 45554 8440 45560 8452
rect 45612 8480 45618 8492
rect 49344 8489 49372 8520
rect 52638 8508 52644 8520
rect 52696 8508 52702 8560
rect 49329 8483 49387 8489
rect 49329 8480 49341 8483
rect 45612 8452 49341 8480
rect 45612 8440 45618 8452
rect 49329 8449 49341 8452
rect 49375 8449 49387 8483
rect 49329 8443 49387 8449
rect 49596 8483 49654 8489
rect 49596 8449 49608 8483
rect 49642 8480 49654 8483
rect 50154 8480 50160 8492
rect 49642 8452 50160 8480
rect 49642 8449 49654 8452
rect 49596 8443 49654 8449
rect 50154 8440 50160 8452
rect 50212 8440 50218 8492
rect 53101 8483 53159 8489
rect 53101 8449 53113 8483
rect 53147 8480 53159 8483
rect 53282 8480 53288 8492
rect 53147 8452 53288 8480
rect 53147 8449 53159 8452
rect 53101 8443 53159 8449
rect 53282 8440 53288 8452
rect 53340 8440 53346 8492
rect 42889 8415 42947 8421
rect 42889 8381 42901 8415
rect 42935 8381 42947 8415
rect 42889 8375 42947 8381
rect 42981 8415 43039 8421
rect 42981 8381 42993 8415
rect 43027 8381 43039 8415
rect 53006 8412 53012 8424
rect 52967 8384 53012 8412
rect 42981 8375 43039 8381
rect 40184 8316 40816 8344
rect 40184 8304 40190 8316
rect 40862 8304 40868 8356
rect 40920 8344 40926 8356
rect 41414 8344 41420 8356
rect 40920 8316 41420 8344
rect 40920 8304 40926 8316
rect 41414 8304 41420 8316
rect 41472 8304 41478 8356
rect 42904 8344 42932 8375
rect 53006 8372 53012 8384
rect 53064 8372 53070 8424
rect 43806 8344 43812 8356
rect 42904 8316 43812 8344
rect 43806 8304 43812 8316
rect 43864 8304 43870 8356
rect 46845 8347 46903 8353
rect 46845 8313 46857 8347
rect 46891 8344 46903 8347
rect 46934 8344 46940 8356
rect 46891 8316 46940 8344
rect 46891 8313 46903 8316
rect 46845 8307 46903 8313
rect 46934 8304 46940 8316
rect 46992 8344 46998 8356
rect 47762 8344 47768 8356
rect 46992 8316 47768 8344
rect 46992 8304 46998 8316
rect 47762 8304 47768 8316
rect 47820 8304 47826 8356
rect 34146 8276 34152 8288
rect 33888 8248 34152 8276
rect 34146 8236 34152 8248
rect 34204 8236 34210 8288
rect 34238 8236 34244 8288
rect 34296 8276 34302 8288
rect 35253 8279 35311 8285
rect 35253 8276 35265 8279
rect 34296 8248 35265 8276
rect 34296 8236 34302 8248
rect 35253 8245 35265 8248
rect 35299 8245 35311 8279
rect 35253 8239 35311 8245
rect 36170 8236 36176 8288
rect 36228 8276 36234 8288
rect 36265 8279 36323 8285
rect 36265 8276 36277 8279
rect 36228 8248 36277 8276
rect 36228 8236 36234 8248
rect 36265 8245 36277 8248
rect 36311 8245 36323 8279
rect 36265 8239 36323 8245
rect 36354 8236 36360 8288
rect 36412 8276 36418 8288
rect 37277 8279 37335 8285
rect 37277 8276 37289 8279
rect 36412 8248 37289 8276
rect 36412 8236 36418 8248
rect 37277 8245 37289 8248
rect 37323 8245 37335 8279
rect 37277 8239 37335 8245
rect 53006 8236 53012 8288
rect 53064 8276 53070 8288
rect 53469 8279 53527 8285
rect 53469 8276 53481 8279
rect 53064 8248 53481 8276
rect 53064 8236 53070 8248
rect 53469 8245 53481 8248
rect 53515 8245 53527 8279
rect 53469 8239 53527 8245
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 3234 8072 3240 8084
rect 3195 8044 3240 8072
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 16908 8044 17509 8072
rect 16908 8032 16914 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 17497 8035 17555 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 26053 8075 26111 8081
rect 26053 8072 26065 8075
rect 24627 8044 24707 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 3252 7936 3280 8032
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 6748 7976 13001 8004
rect 3252 7908 4200 7936
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 1946 7868 1952 7880
rect 1903 7840 1952 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 4172 7877 4200 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4614 7868 4620 7880
rect 4295 7840 4620 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 2124 7803 2182 7809
rect 2124 7769 2136 7803
rect 2170 7800 2182 7803
rect 3789 7803 3847 7809
rect 3789 7800 3801 7803
rect 2170 7772 3801 7800
rect 2170 7769 2182 7772
rect 2124 7763 2182 7769
rect 3789 7769 3801 7772
rect 3835 7769 3847 7803
rect 3988 7800 4016 7831
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 6748 7877 6776 7976
rect 12989 7973 13001 7976
rect 13035 7973 13047 8007
rect 12989 7967 13047 7973
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 13780 7976 16528 8004
rect 13780 7964 13786 7976
rect 13078 7936 13084 7948
rect 6840 7908 13084 7936
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6840 7800 6868 7908
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 14550 7936 14556 7948
rect 13403 7908 14556 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 15988 7908 16221 7936
rect 15988 7896 15994 7908
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7466 7868 7472 7880
rect 7055 7840 7472 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 9858 7868 9864 7880
rect 9819 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10594 7868 10600 7880
rect 10275 7840 10600 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10594 7828 10600 7840
rect 10652 7868 10658 7880
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 10652 7840 10793 7868
rect 10652 7828 10658 7840
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11480 7840 11621 7868
rect 11480 7828 11486 7840
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 13170 7868 13176 7880
rect 13131 7840 13176 7868
rect 11793 7831 11851 7837
rect 3988 7772 6868 7800
rect 3789 7763 3847 7769
rect 9950 7760 9956 7812
rect 10008 7800 10014 7812
rect 11808 7800 11836 7831
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 13449 7871 13507 7877
rect 13320 7840 13365 7868
rect 13320 7828 13326 7840
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 14090 7868 14096 7880
rect 14051 7840 14096 7868
rect 13449 7831 13507 7837
rect 10008 7772 11836 7800
rect 13464 7800 13492 7831
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 16500 7877 16528 7976
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 24679 8004 24707 8044
rect 24877 8044 26065 8072
rect 24877 8004 24905 8044
rect 26053 8041 26065 8044
rect 26099 8041 26111 8075
rect 26053 8035 26111 8041
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 28629 8075 28687 8081
rect 28629 8072 28641 8075
rect 28132 8044 28641 8072
rect 28132 8032 28138 8044
rect 28629 8041 28641 8044
rect 28675 8041 28687 8075
rect 28629 8035 28687 8041
rect 28718 8032 28724 8084
rect 28776 8072 28782 8084
rect 33042 8072 33048 8084
rect 28776 8044 31754 8072
rect 33003 8044 33048 8072
rect 28776 8032 28782 8044
rect 30282 8004 30288 8016
rect 17276 7976 17816 8004
rect 24679 7976 24905 8004
rect 24964 7976 30288 8004
rect 17276 7964 17282 7976
rect 17678 7936 17684 7948
rect 17639 7908 17684 7936
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17788 7945 17816 7976
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 18414 7936 18420 7948
rect 18003 7908 18420 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7936 21603 7939
rect 24489 7939 24547 7945
rect 24489 7936 24501 7939
rect 21591 7908 24501 7936
rect 21591 7905 21603 7908
rect 21545 7899 21603 7905
rect 24489 7905 24501 7908
rect 24535 7936 24547 7939
rect 24964 7936 24992 7976
rect 30282 7964 30288 7976
rect 30340 7964 30346 8016
rect 31726 8004 31754 8044
rect 33042 8032 33048 8044
rect 33100 8032 33106 8084
rect 33502 8032 33508 8084
rect 33560 8072 33566 8084
rect 36449 8075 36507 8081
rect 36449 8072 36461 8075
rect 33560 8044 36461 8072
rect 33560 8032 33566 8044
rect 36449 8041 36461 8044
rect 36495 8072 36507 8075
rect 40586 8072 40592 8084
rect 36495 8044 40592 8072
rect 36495 8041 36507 8044
rect 36449 8035 36507 8041
rect 40586 8032 40592 8044
rect 40644 8032 40650 8084
rect 42242 8072 42248 8084
rect 42203 8044 42248 8072
rect 42242 8032 42248 8044
rect 42300 8032 42306 8084
rect 50154 8072 50160 8084
rect 50115 8044 50160 8072
rect 50154 8032 50160 8044
rect 50212 8032 50218 8084
rect 53282 8032 53288 8084
rect 53340 8072 53346 8084
rect 54021 8075 54079 8081
rect 54021 8072 54033 8075
rect 53340 8044 54033 8072
rect 53340 8032 53346 8044
rect 54021 8041 54033 8044
rect 54067 8041 54079 8075
rect 54021 8035 54079 8041
rect 49510 8004 49516 8016
rect 31726 7976 49516 8004
rect 49510 7964 49516 7976
rect 49568 8004 49574 8016
rect 50525 8007 50583 8013
rect 50525 8004 50537 8007
rect 49568 7976 50537 8004
rect 49568 7964 49574 7976
rect 50525 7973 50537 7976
rect 50571 8004 50583 8007
rect 50706 8004 50712 8016
rect 50571 7976 50712 8004
rect 50571 7973 50583 7976
rect 50525 7967 50583 7973
rect 50706 7964 50712 7976
rect 50764 7964 50770 8016
rect 27522 7936 27528 7948
rect 24535 7908 24992 7936
rect 26068 7908 27528 7936
rect 24535 7905 24547 7908
rect 24489 7899 24547 7905
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 14240 7840 14381 7868
rect 14240 7828 14246 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7868 16543 7871
rect 16666 7868 16672 7880
rect 16531 7840 16672 7868
rect 16531 7837 16543 7840
rect 16485 7831 16543 7837
rect 16666 7828 16672 7840
rect 16724 7868 16730 7880
rect 17126 7868 17132 7880
rect 16724 7840 17132 7868
rect 16724 7828 16730 7840
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 16114 7800 16120 7812
rect 13464 7772 16120 7800
rect 10008 7760 10014 7772
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16206 7760 16212 7812
rect 16264 7800 16270 7812
rect 17310 7800 17316 7812
rect 16264 7772 17316 7800
rect 16264 7760 16270 7772
rect 17310 7760 17316 7772
rect 17368 7760 17374 7812
rect 6549 7735 6607 7741
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 6638 7732 6644 7744
rect 6595 7704 6644 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 11054 7732 11060 7744
rect 6972 7704 7017 7732
rect 11015 7704 11060 7732
rect 6972 7692 6978 7704
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11572 7704 11713 7732
rect 11572 7692 11578 7704
rect 11701 7701 11713 7704
rect 11747 7701 11759 7735
rect 11701 7695 11759 7701
rect 17770 7692 17776 7744
rect 17828 7732 17834 7744
rect 17880 7732 17908 7831
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19392 7840 19625 7868
rect 19392 7828 19398 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 19880 7803 19938 7809
rect 19880 7769 19892 7803
rect 19926 7800 19938 7803
rect 20806 7800 20812 7812
rect 19926 7772 20812 7800
rect 19926 7769 19938 7772
rect 19880 7763 19938 7769
rect 20806 7760 20812 7772
rect 20864 7760 20870 7812
rect 21468 7800 21496 7831
rect 22738 7828 22744 7880
rect 22796 7868 22802 7880
rect 26068 7877 26096 7908
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 27798 7896 27804 7948
rect 27856 7936 27862 7948
rect 33594 7936 33600 7948
rect 27856 7908 28856 7936
rect 33555 7908 33600 7936
rect 27856 7896 27862 7908
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 22796 7840 24409 7868
rect 22796 7828 22802 7840
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 26053 7871 26111 7877
rect 26053 7837 26065 7871
rect 26099 7837 26111 7871
rect 26053 7831 26111 7837
rect 26237 7871 26295 7877
rect 26237 7837 26249 7871
rect 26283 7837 26295 7871
rect 26878 7868 26884 7880
rect 26839 7840 26884 7868
rect 26237 7831 26295 7837
rect 22186 7800 22192 7812
rect 21468 7772 22192 7800
rect 22186 7760 22192 7772
rect 22244 7760 22250 7812
rect 25130 7760 25136 7812
rect 25188 7800 25194 7812
rect 26252 7800 26280 7831
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 27154 7868 27160 7880
rect 27115 7840 27160 7868
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7868 28043 7871
rect 28166 7868 28172 7880
rect 28031 7840 28172 7868
rect 28031 7837 28043 7840
rect 27985 7831 28043 7837
rect 28166 7828 28172 7840
rect 28224 7828 28230 7880
rect 28626 7868 28632 7880
rect 28587 7840 28632 7868
rect 28626 7828 28632 7840
rect 28684 7828 28690 7880
rect 28828 7877 28856 7908
rect 33594 7896 33600 7908
rect 33652 7936 33658 7948
rect 38749 7939 38807 7945
rect 38749 7936 38761 7939
rect 33652 7908 38761 7936
rect 33652 7896 33658 7908
rect 38749 7905 38761 7908
rect 38795 7936 38807 7939
rect 39114 7936 39120 7948
rect 38795 7908 39120 7936
rect 38795 7905 38807 7908
rect 38749 7899 38807 7905
rect 39114 7896 39120 7908
rect 39172 7896 39178 7948
rect 40034 7896 40040 7948
rect 40092 7936 40098 7948
rect 40678 7936 40684 7948
rect 40092 7908 40684 7936
rect 40092 7896 40098 7908
rect 40678 7896 40684 7908
rect 40736 7896 40742 7948
rect 42702 7896 42708 7948
rect 42760 7936 42766 7948
rect 42797 7939 42855 7945
rect 42797 7936 42809 7939
rect 42760 7908 42809 7936
rect 42760 7896 42766 7908
rect 42797 7905 42809 7908
rect 42843 7905 42855 7939
rect 50614 7936 50620 7948
rect 50575 7908 50620 7936
rect 42797 7899 42855 7905
rect 50614 7896 50620 7908
rect 50672 7896 50678 7948
rect 52638 7936 52644 7948
rect 52599 7908 52644 7936
rect 52638 7896 52644 7908
rect 52696 7896 52702 7948
rect 28813 7871 28871 7877
rect 28813 7837 28825 7871
rect 28859 7837 28871 7871
rect 28813 7831 28871 7837
rect 30466 7828 30472 7880
rect 30524 7868 30530 7880
rect 36170 7868 36176 7880
rect 30524 7840 36176 7868
rect 30524 7828 30530 7840
rect 36170 7828 36176 7840
rect 36228 7828 36234 7880
rect 36265 7871 36323 7877
rect 36265 7837 36277 7871
rect 36311 7868 36323 7871
rect 36354 7868 36360 7880
rect 36311 7840 36360 7868
rect 36311 7837 36323 7840
rect 36265 7831 36323 7837
rect 36354 7828 36360 7840
rect 36412 7828 36418 7880
rect 38378 7828 38384 7880
rect 38436 7868 38442 7880
rect 38565 7871 38623 7877
rect 38565 7868 38577 7871
rect 38436 7840 38577 7868
rect 38436 7828 38442 7840
rect 38565 7837 38577 7840
rect 38611 7837 38623 7871
rect 38565 7831 38623 7837
rect 50246 7828 50252 7880
rect 50304 7868 50310 7880
rect 50341 7871 50399 7877
rect 50341 7868 50353 7871
rect 50304 7840 50353 7868
rect 50304 7828 50310 7840
rect 50341 7837 50353 7840
rect 50387 7837 50399 7871
rect 50341 7831 50399 7837
rect 27617 7803 27675 7809
rect 27617 7800 27629 7803
rect 25188 7772 27629 7800
rect 25188 7760 25194 7772
rect 27617 7769 27629 7772
rect 27663 7769 27675 7803
rect 27617 7763 27675 7769
rect 27893 7803 27951 7809
rect 27893 7769 27905 7803
rect 27939 7800 27951 7803
rect 29546 7800 29552 7812
rect 27939 7772 29552 7800
rect 27939 7769 27951 7772
rect 27893 7763 27951 7769
rect 29546 7760 29552 7772
rect 29604 7760 29610 7812
rect 33226 7760 33232 7812
rect 33284 7800 33290 7812
rect 33505 7803 33563 7809
rect 33505 7800 33517 7803
rect 33284 7772 33517 7800
rect 33284 7760 33290 7772
rect 33505 7769 33517 7772
rect 33551 7769 33563 7803
rect 42610 7800 42616 7812
rect 42523 7772 42616 7800
rect 33505 7763 33563 7769
rect 42610 7760 42616 7772
rect 42668 7800 42674 7812
rect 45186 7800 45192 7812
rect 42668 7772 45192 7800
rect 42668 7760 42674 7772
rect 45186 7760 45192 7772
rect 45244 7760 45250 7812
rect 52908 7803 52966 7809
rect 52908 7769 52920 7803
rect 52954 7800 52966 7803
rect 53098 7800 53104 7812
rect 52954 7772 53104 7800
rect 52954 7769 52966 7772
rect 52908 7763 52966 7769
rect 53098 7760 53104 7772
rect 53156 7760 53162 7812
rect 20990 7732 20996 7744
rect 17828 7704 17908 7732
rect 20951 7704 20996 7732
rect 17828 7692 17834 7704
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 21818 7732 21824 7744
rect 21779 7704 21824 7732
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 23842 7692 23848 7744
rect 23900 7732 23906 7744
rect 24765 7735 24823 7741
rect 24765 7732 24777 7735
rect 23900 7704 24777 7732
rect 23900 7692 23906 7704
rect 24765 7701 24777 7704
rect 24811 7701 24823 7735
rect 26694 7732 26700 7744
rect 26655 7704 26700 7732
rect 24765 7695 24823 7701
rect 26694 7692 26700 7704
rect 26752 7692 26758 7744
rect 27062 7732 27068 7744
rect 27023 7704 27068 7732
rect 27062 7692 27068 7704
rect 27120 7692 27126 7744
rect 27798 7732 27804 7744
rect 27759 7704 27804 7732
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 28166 7732 28172 7744
rect 28127 7704 28172 7732
rect 28166 7692 28172 7704
rect 28224 7692 28230 7744
rect 33413 7735 33471 7741
rect 33413 7701 33425 7735
rect 33459 7732 33471 7735
rect 34330 7732 34336 7744
rect 33459 7704 34336 7732
rect 33459 7701 33471 7704
rect 33413 7695 33471 7701
rect 34330 7692 34336 7704
rect 34388 7692 34394 7744
rect 42705 7735 42763 7741
rect 42705 7701 42717 7735
rect 42751 7732 42763 7735
rect 42794 7732 42800 7744
rect 42751 7704 42800 7732
rect 42751 7701 42763 7704
rect 42705 7695 42763 7701
rect 42794 7692 42800 7704
rect 42852 7732 42858 7744
rect 43898 7732 43904 7744
rect 42852 7704 43904 7732
rect 42852 7692 42858 7704
rect 43898 7692 43904 7704
rect 43956 7692 43962 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 12710 7528 12716 7540
rect 2823 7500 12716 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13725 7531 13783 7537
rect 13725 7528 13737 7531
rect 13228 7500 13737 7528
rect 13228 7488 13234 7500
rect 13725 7497 13737 7500
rect 13771 7497 13783 7531
rect 13725 7491 13783 7497
rect 16850 7488 16856 7540
rect 16908 7488 16914 7540
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 35437 7531 35495 7537
rect 35437 7528 35449 7531
rect 22066 7500 35449 7528
rect 6914 7460 6920 7472
rect 1412 7432 6920 7460
rect 1412 7401 1440 7432
rect 6914 7420 6920 7432
rect 6972 7460 6978 7472
rect 14274 7460 14280 7472
rect 6972 7432 7788 7460
rect 6972 7420 6978 7432
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 2314 7392 2320 7404
rect 2275 7364 2320 7392
rect 1397 7355 1455 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 2958 7392 2964 7404
rect 2919 7364 2964 7392
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 6362 7392 6368 7404
rect 6323 7364 6368 7392
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6638 7401 6644 7404
rect 6632 7392 6644 7401
rect 6599 7364 6644 7392
rect 6632 7355 6644 7364
rect 6638 7352 6644 7355
rect 6696 7352 6702 7404
rect 2133 7259 2191 7265
rect 2133 7225 2145 7259
rect 2179 7256 2191 7259
rect 3234 7256 3240 7268
rect 2179 7228 3240 7256
rect 2179 7225 2191 7228
rect 2133 7219 2191 7225
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 7760 7265 7788 7432
rect 14016 7432 14280 7460
rect 9674 7401 9680 7404
rect 9668 7355 9680 7401
rect 9732 7392 9738 7404
rect 13906 7392 13912 7404
rect 9732 7364 9768 7392
rect 13867 7364 13912 7392
rect 9674 7352 9680 7355
rect 9732 7352 9738 7364
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14016 7401 14044 7432
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 16868 7460 16896 7488
rect 16945 7463 17003 7469
rect 16945 7460 16957 7463
rect 16868 7432 16957 7460
rect 16945 7429 16957 7432
rect 16991 7429 17003 7463
rect 16945 7423 17003 7429
rect 17037 7463 17095 7469
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 19242 7460 19248 7472
rect 17083 7432 19248 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14458 7392 14464 7404
rect 14139 7364 14464 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 15289 7395 15347 7401
rect 15289 7392 15301 7395
rect 15252 7364 15301 7392
rect 15252 7352 15258 7364
rect 15289 7361 15301 7364
rect 15335 7361 15347 7395
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 15289 7355 15347 7361
rect 16132 7364 16681 7392
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7324 14243 7327
rect 14642 7324 14648 7336
rect 14231 7296 14648 7324
rect 14231 7293 14243 7296
rect 14185 7287 14243 7293
rect 7745 7259 7803 7265
rect 7745 7225 7757 7259
rect 7791 7225 7803 7259
rect 7745 7219 7803 7225
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6362 7188 6368 7200
rect 6144 7160 6368 7188
rect 6144 7148 6150 7160
rect 6362 7148 6368 7160
rect 6420 7188 6426 7200
rect 9416 7188 9444 7287
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 10781 7259 10839 7265
rect 10781 7225 10793 7259
rect 10827 7256 10839 7259
rect 11422 7256 11428 7268
rect 10827 7228 11428 7256
rect 10827 7225 10839 7228
rect 10781 7219 10839 7225
rect 11422 7216 11428 7228
rect 11480 7216 11486 7268
rect 14090 7216 14096 7268
rect 14148 7256 14154 7268
rect 15580 7256 15608 7287
rect 16132 7268 16160 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16817 7395 16875 7401
rect 16817 7361 16829 7395
rect 16863 7361 16875 7395
rect 16817 7355 16875 7361
rect 16832 7324 16860 7355
rect 17126 7352 17132 7404
rect 17184 7401 17190 7404
rect 17184 7392 17192 7401
rect 17678 7392 17684 7404
rect 17184 7364 17684 7392
rect 17184 7355 17192 7364
rect 17184 7352 17190 7355
rect 17678 7352 17684 7364
rect 17736 7352 17742 7404
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 19886 7324 19892 7336
rect 16832 7296 19892 7324
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 20548 7324 20576 7355
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20680 7364 20725 7392
rect 20680 7352 20686 7364
rect 20714 7324 20720 7336
rect 20548 7296 20720 7324
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7324 20867 7327
rect 21818 7324 21824 7336
rect 20855 7296 21824 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 21818 7284 21824 7296
rect 21876 7284 21882 7336
rect 16114 7256 16120 7268
rect 14148 7228 16120 7256
rect 14148 7216 14154 7228
rect 16114 7216 16120 7228
rect 16172 7216 16178 7268
rect 22066 7256 22094 7500
rect 35437 7497 35449 7500
rect 35483 7528 35495 7531
rect 36015 7531 36073 7537
rect 35483 7500 35848 7528
rect 35483 7497 35495 7500
rect 35437 7491 35495 7497
rect 22480 7432 22876 7460
rect 22480 7404 22508 7432
rect 22462 7392 22468 7404
rect 22375 7364 22468 7392
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 22738 7392 22744 7404
rect 22699 7364 22744 7392
rect 22738 7352 22744 7364
rect 22796 7352 22802 7404
rect 22848 7392 22876 7432
rect 23750 7420 23756 7472
rect 23808 7460 23814 7472
rect 23998 7463 24056 7469
rect 23998 7460 24010 7463
rect 23808 7432 24010 7460
rect 23808 7420 23814 7432
rect 23998 7429 24010 7432
rect 24044 7429 24056 7463
rect 23998 7423 24056 7429
rect 26694 7420 26700 7472
rect 26752 7460 26758 7472
rect 27218 7463 27276 7469
rect 27218 7460 27230 7463
rect 26752 7432 27230 7460
rect 26752 7420 26758 7432
rect 27218 7429 27230 7432
rect 27264 7429 27276 7463
rect 27218 7423 27276 7429
rect 27706 7420 27712 7472
rect 27764 7460 27770 7472
rect 28626 7460 28632 7472
rect 27764 7432 28632 7460
rect 27764 7420 27770 7432
rect 28626 7420 28632 7432
rect 28684 7420 28690 7472
rect 32493 7463 32551 7469
rect 32493 7429 32505 7463
rect 32539 7460 32551 7463
rect 32858 7460 32864 7472
rect 32539 7432 32864 7460
rect 32539 7429 32551 7432
rect 32493 7423 32551 7429
rect 32858 7420 32864 7432
rect 32916 7420 32922 7472
rect 35820 7469 35848 7500
rect 36015 7497 36027 7531
rect 36061 7528 36073 7531
rect 36354 7528 36360 7540
rect 36061 7500 36360 7528
rect 36061 7497 36073 7500
rect 36015 7491 36073 7497
rect 36354 7488 36360 7500
rect 36412 7488 36418 7540
rect 36538 7488 36544 7540
rect 36596 7528 36602 7540
rect 36998 7528 37004 7540
rect 36596 7500 37004 7528
rect 36596 7488 36602 7500
rect 36998 7488 37004 7500
rect 37056 7488 37062 7540
rect 53098 7528 53104 7540
rect 53059 7500 53104 7528
rect 53098 7488 53104 7500
rect 53156 7488 53162 7540
rect 35805 7463 35863 7469
rect 35805 7429 35817 7463
rect 35851 7429 35863 7463
rect 35805 7423 35863 7429
rect 36446 7420 36452 7472
rect 36504 7460 36510 7472
rect 37090 7460 37096 7472
rect 36504 7432 37096 7460
rect 36504 7420 36510 7432
rect 37090 7420 37096 7432
rect 37148 7420 37154 7472
rect 37458 7420 37464 7472
rect 37516 7460 37522 7472
rect 37737 7463 37795 7469
rect 37737 7460 37749 7463
rect 37516 7432 37749 7460
rect 37516 7420 37522 7432
rect 37737 7429 37749 7432
rect 37783 7429 37795 7463
rect 37737 7423 37795 7429
rect 40678 7420 40684 7472
rect 40736 7460 40742 7472
rect 43962 7463 44020 7469
rect 43962 7460 43974 7463
rect 40736 7432 43974 7460
rect 40736 7420 40742 7432
rect 43962 7429 43974 7432
rect 44008 7429 44020 7463
rect 43962 7423 44020 7429
rect 52914 7420 52920 7472
rect 52972 7460 52978 7472
rect 52972 7432 53236 7460
rect 52972 7420 52978 7432
rect 28166 7392 28172 7404
rect 22848 7364 28172 7392
rect 28166 7352 28172 7364
rect 28224 7352 28230 7404
rect 32306 7392 32312 7404
rect 32267 7364 32312 7392
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 32631 7395 32689 7401
rect 32456 7364 32501 7392
rect 32456 7352 32462 7364
rect 32631 7361 32643 7395
rect 32677 7361 32689 7395
rect 32631 7355 32689 7361
rect 21836 7228 22094 7256
rect 9582 7188 9588 7200
rect 6420 7160 9588 7188
rect 6420 7148 6426 7160
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 21836 7188 21864 7228
rect 12584 7160 21864 7188
rect 12584 7148 12590 7160
rect 21910 7148 21916 7200
rect 21968 7188 21974 7200
rect 22756 7188 22784 7352
rect 23474 7284 23480 7336
rect 23532 7324 23538 7336
rect 23753 7327 23811 7333
rect 23753 7324 23765 7327
rect 23532 7296 23765 7324
rect 23532 7284 23538 7296
rect 23753 7293 23765 7296
rect 23799 7293 23811 7327
rect 23753 7287 23811 7293
rect 26786 7284 26792 7336
rect 26844 7324 26850 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26844 7296 26985 7324
rect 26844 7284 26850 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 30926 7284 30932 7336
rect 30984 7324 30990 7336
rect 32490 7324 32496 7336
rect 30984 7296 32496 7324
rect 30984 7284 30990 7296
rect 32490 7284 32496 7296
rect 32548 7324 32554 7336
rect 32646 7324 32674 7355
rect 33134 7352 33140 7404
rect 33192 7392 33198 7404
rect 33597 7395 33655 7401
rect 33597 7392 33609 7395
rect 33192 7364 33609 7392
rect 33192 7352 33198 7364
rect 33597 7361 33609 7364
rect 33643 7361 33655 7395
rect 33597 7355 33655 7361
rect 35434 7352 35440 7404
rect 35492 7392 35498 7404
rect 37476 7392 37504 7420
rect 35492 7364 37504 7392
rect 35492 7352 35498 7364
rect 38378 7352 38384 7404
rect 38436 7392 38442 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 38436 7364 38577 7392
rect 38436 7352 38442 7364
rect 38565 7361 38577 7364
rect 38611 7361 38623 7395
rect 43714 7392 43720 7404
rect 43675 7364 43720 7392
rect 38565 7355 38623 7361
rect 43714 7352 43720 7364
rect 43772 7352 43778 7404
rect 44542 7352 44548 7404
rect 44600 7392 44606 7404
rect 45278 7392 45284 7404
rect 44600 7364 45284 7392
rect 44600 7352 44606 7364
rect 45278 7352 45284 7364
rect 45336 7392 45342 7404
rect 46385 7395 46443 7401
rect 46385 7392 46397 7395
rect 45336 7364 46397 7392
rect 45336 7352 45342 7364
rect 46385 7361 46397 7364
rect 46431 7392 46443 7395
rect 47302 7392 47308 7404
rect 46431 7364 47308 7392
rect 46431 7361 46443 7364
rect 46385 7355 46443 7361
rect 47302 7352 47308 7364
rect 47360 7352 47366 7404
rect 53006 7392 53012 7404
rect 52967 7364 53012 7392
rect 53006 7352 53012 7364
rect 53064 7352 53070 7404
rect 53208 7401 53236 7432
rect 53193 7395 53251 7401
rect 53193 7361 53205 7395
rect 53239 7361 53251 7395
rect 53193 7355 53251 7361
rect 32548 7296 32674 7324
rect 32769 7327 32827 7333
rect 32548 7284 32554 7296
rect 32769 7293 32781 7327
rect 32815 7293 32827 7327
rect 32769 7287 32827 7293
rect 46661 7327 46719 7333
rect 46661 7293 46673 7327
rect 46707 7324 46719 7327
rect 46934 7324 46940 7336
rect 46707 7296 46940 7324
rect 46707 7293 46719 7296
rect 46661 7287 46719 7293
rect 32784 7256 32812 7287
rect 46934 7284 46940 7296
rect 46992 7284 46998 7336
rect 24688 7228 25268 7256
rect 21968 7160 22784 7188
rect 21968 7148 21974 7160
rect 22922 7148 22928 7200
rect 22980 7188 22986 7200
rect 24688 7188 24716 7228
rect 25130 7188 25136 7200
rect 22980 7160 24716 7188
rect 25091 7160 25136 7188
rect 22980 7148 22986 7160
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 25240 7188 25268 7228
rect 27908 7228 32812 7256
rect 33781 7259 33839 7265
rect 27908 7188 27936 7228
rect 33781 7225 33793 7259
rect 33827 7256 33839 7259
rect 35342 7256 35348 7268
rect 33827 7228 35348 7256
rect 33827 7225 33839 7228
rect 33781 7219 33839 7225
rect 25240 7160 27936 7188
rect 27982 7148 27988 7200
rect 28040 7188 28046 7200
rect 28353 7191 28411 7197
rect 28353 7188 28365 7191
rect 28040 7160 28365 7188
rect 28040 7148 28046 7160
rect 28353 7157 28365 7160
rect 28399 7157 28411 7191
rect 32122 7188 32128 7200
rect 32083 7160 32128 7188
rect 28353 7151 28411 7157
rect 32122 7148 32128 7160
rect 32180 7148 32186 7200
rect 32398 7148 32404 7200
rect 32456 7188 32462 7200
rect 33318 7188 33324 7200
rect 32456 7160 33324 7188
rect 32456 7148 32462 7160
rect 33318 7148 33324 7160
rect 33376 7188 33382 7200
rect 33796 7188 33824 7219
rect 35342 7216 35348 7228
rect 35400 7216 35406 7268
rect 36998 7216 37004 7268
rect 37056 7256 37062 7268
rect 38749 7259 38807 7265
rect 38749 7256 38761 7259
rect 37056 7228 38761 7256
rect 37056 7216 37062 7228
rect 38749 7225 38761 7228
rect 38795 7256 38807 7259
rect 42702 7256 42708 7268
rect 38795 7228 42708 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 42702 7216 42708 7228
rect 42760 7216 42766 7268
rect 35986 7188 35992 7200
rect 33376 7160 33824 7188
rect 35947 7160 35992 7188
rect 33376 7148 33382 7160
rect 35986 7148 35992 7160
rect 36044 7148 36050 7200
rect 36170 7188 36176 7200
rect 36131 7160 36176 7188
rect 36170 7148 36176 7160
rect 36228 7148 36234 7200
rect 37826 7188 37832 7200
rect 37787 7160 37832 7188
rect 37826 7148 37832 7160
rect 37884 7148 37890 7200
rect 45097 7191 45155 7197
rect 45097 7157 45109 7191
rect 45143 7188 45155 7191
rect 45186 7188 45192 7200
rect 45143 7160 45192 7188
rect 45143 7157 45155 7160
rect 45097 7151 45155 7157
rect 45186 7148 45192 7160
rect 45244 7148 45250 7200
rect 46198 7188 46204 7200
rect 46159 7160 46204 7188
rect 46198 7148 46204 7160
rect 46256 7148 46262 7200
rect 46566 7188 46572 7200
rect 46527 7160 46572 7188
rect 46566 7148 46572 7160
rect 46624 7148 46630 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 9732 6956 9781 6984
rect 9732 6944 9738 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13320 6956 13553 6984
rect 13320 6944 13326 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14642 6984 14648 6996
rect 13780 6956 14648 6984
rect 13780 6944 13786 6956
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 16114 6944 16120 6996
rect 16172 6984 16178 6996
rect 16172 6956 17264 6984
rect 16172 6944 16178 6956
rect 2038 6876 2044 6928
rect 2096 6916 2102 6928
rect 3786 6916 3792 6928
rect 2096 6888 3792 6916
rect 2096 6876 2102 6888
rect 3786 6876 3792 6888
rect 3844 6876 3850 6928
rect 8018 6876 8024 6928
rect 8076 6916 8082 6928
rect 9950 6916 9956 6928
rect 8076 6888 9956 6916
rect 8076 6876 8082 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 16206 6876 16212 6928
rect 16264 6876 16270 6928
rect 16850 6916 16856 6928
rect 16408 6888 16856 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 9674 6848 9680 6860
rect 1719 6820 3924 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 2832 6752 3157 6780
rect 2832 6740 2838 6752
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3786 6780 3792 6792
rect 3747 6752 3792 6780
rect 3145 6743 3203 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3896 6780 3924 6820
rect 4816 6820 9680 6848
rect 4816 6780 4844 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9968 6848 9996 6876
rect 14918 6848 14924 6860
rect 9784 6820 9996 6848
rect 12912 6820 14044 6848
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 3896 6752 4844 6780
rect 5184 6752 6469 6780
rect 4034 6715 4092 6721
rect 4034 6712 4046 6715
rect 2976 6684 4046 6712
rect 2976 6653 3004 6684
rect 4034 6681 4046 6684
rect 4080 6681 4092 6715
rect 4034 6675 4092 6681
rect 5184 6656 5212 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7098 6780 7104 6792
rect 6779 6752 7104 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 6656 6712 6684 6743
rect 7098 6740 7104 6752
rect 7156 6780 7162 6792
rect 7466 6780 7472 6792
rect 7156 6752 7472 6780
rect 7156 6740 7162 6752
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 9784 6789 9812 6820
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6780 10011 6783
rect 11054 6780 11060 6792
rect 9999 6752 11060 6780
rect 9999 6749 10011 6752
rect 9953 6743 10011 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 12912 6789 12940 6820
rect 13078 6789 13084 6792
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13045 6783 13084 6789
rect 13045 6749 13057 6783
rect 13045 6743 13084 6749
rect 13078 6740 13084 6743
rect 13136 6740 13142 6792
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13403 6783 13461 6789
rect 13403 6749 13415 6783
rect 13449 6780 13461 6783
rect 13722 6780 13728 6792
rect 13449 6752 13728 6780
rect 13449 6749 13461 6752
rect 13403 6743 13461 6749
rect 7834 6712 7840 6724
rect 6656 6684 7840 6712
rect 7834 6672 7840 6684
rect 7892 6672 7898 6724
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6613 3019 6647
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 2961 6607 3019 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 9950 6644 9956 6656
rect 7156 6616 9956 6644
rect 7156 6604 7162 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 13188 6644 13216 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 14016 6780 14044 6820
rect 14476 6820 14924 6848
rect 14090 6780 14096 6792
rect 14148 6789 14154 6792
rect 14003 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6743 14158 6789
rect 14186 6783 14244 6789
rect 14186 6749 14198 6783
rect 14232 6780 14244 6783
rect 14274 6780 14280 6792
rect 14232 6752 14280 6780
rect 14232 6749 14244 6752
rect 14186 6743 14244 6749
rect 14148 6740 14154 6743
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14476 6789 14504 6820
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 14642 6789 14648 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14599 6783 14648 6789
rect 14599 6749 14611 6783
rect 14645 6749 14648 6783
rect 14599 6743 14648 6749
rect 14642 6740 14648 6743
rect 14700 6740 14706 6792
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16224 6789 16252 6876
rect 16210 6783 16268 6789
rect 16210 6749 16222 6783
rect 16256 6749 16268 6783
rect 16210 6743 16268 6749
rect 13262 6672 13268 6724
rect 13320 6712 13326 6724
rect 16408 6721 16436 6888
rect 16832 6876 16856 6888
rect 16908 6916 16914 6928
rect 16908 6888 16965 6916
rect 16908 6876 16914 6888
rect 16666 6789 16672 6792
rect 16623 6783 16672 6789
rect 16623 6749 16635 6783
rect 16669 6749 16672 6783
rect 16623 6743 16672 6749
rect 16666 6740 16672 6743
rect 16724 6740 16730 6792
rect 14369 6715 14427 6721
rect 13320 6684 13365 6712
rect 13320 6672 13326 6684
rect 14369 6681 14381 6715
rect 14415 6681 14427 6715
rect 16393 6715 16451 6721
rect 16393 6712 16405 6715
rect 14369 6675 14427 6681
rect 14568 6684 16405 6712
rect 14182 6644 14188 6656
rect 13188 6616 14188 6644
rect 14182 6604 14188 6616
rect 14240 6644 14246 6656
rect 14384 6644 14412 6675
rect 14568 6644 14596 6684
rect 16393 6681 16405 6684
rect 16439 6681 16451 6715
rect 16393 6675 16451 6681
rect 16485 6715 16543 6721
rect 16485 6681 16497 6715
rect 16531 6712 16543 6715
rect 16832 6712 16860 6876
rect 17236 6789 17264 6956
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 20349 6987 20407 6993
rect 20349 6984 20361 6987
rect 19484 6956 20361 6984
rect 19484 6944 19490 6956
rect 20349 6953 20361 6956
rect 20395 6953 20407 6987
rect 21542 6984 21548 6996
rect 21503 6956 21548 6984
rect 20349 6947 20407 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 21634 6944 21640 6996
rect 21692 6984 21698 6996
rect 25130 6984 25136 6996
rect 21692 6956 25136 6984
rect 21692 6944 21698 6956
rect 25130 6944 25136 6956
rect 25188 6944 25194 6996
rect 32306 6944 32312 6996
rect 32364 6984 32370 6996
rect 32861 6987 32919 6993
rect 32861 6984 32873 6987
rect 32364 6956 32873 6984
rect 32364 6944 32370 6956
rect 32861 6953 32873 6956
rect 32907 6953 32919 6987
rect 35986 6984 35992 6996
rect 35947 6956 35992 6984
rect 32861 6947 32919 6953
rect 35986 6944 35992 6956
rect 36044 6944 36050 6996
rect 36170 6944 36176 6996
rect 36228 6984 36234 6996
rect 46566 6984 46572 6996
rect 36228 6956 46572 6984
rect 36228 6944 36234 6956
rect 46566 6944 46572 6956
rect 46624 6944 46630 6996
rect 20990 6916 20996 6928
rect 19306 6888 20996 6916
rect 19306 6848 19334 6888
rect 20990 6876 20996 6888
rect 21048 6876 21054 6928
rect 36998 6916 37004 6928
rect 33520 6888 37004 6916
rect 21910 6848 21916 6860
rect 17420 6820 19334 6848
rect 20456 6820 21916 6848
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17420 6780 17448 6820
rect 17368 6752 17448 6780
rect 17368 6740 17374 6752
rect 17678 6740 17684 6792
rect 17736 6789 17742 6792
rect 17736 6780 17744 6789
rect 17736 6752 17781 6780
rect 17736 6743 17744 6752
rect 17736 6740 17742 6743
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 20254 6780 20260 6792
rect 19944 6752 20260 6780
rect 19944 6740 19950 6752
rect 17497 6715 17555 6721
rect 17497 6712 17509 6715
rect 16531 6684 16712 6712
rect 16832 6684 17509 6712
rect 16531 6681 16543 6684
rect 16485 6675 16543 6681
rect 16684 6656 16712 6684
rect 17497 6681 17509 6684
rect 17543 6681 17555 6715
rect 17497 6675 17555 6681
rect 17589 6715 17647 6721
rect 17589 6681 17601 6715
rect 17635 6712 17647 6715
rect 20070 6712 20076 6724
rect 17635 6684 20076 6712
rect 17635 6681 17647 6684
rect 17589 6675 17647 6681
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20180 6721 20208 6752
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6681 20223 6715
rect 20165 6675 20223 6681
rect 20370 6715 20428 6721
rect 20370 6681 20382 6715
rect 20416 6712 20428 6715
rect 20456 6712 20484 6820
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22186 6848 22192 6860
rect 22147 6820 22192 6848
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 26050 6808 26056 6860
rect 26108 6848 26114 6860
rect 30926 6848 30932 6860
rect 26108 6820 30932 6848
rect 26108 6808 26114 6820
rect 30926 6808 30932 6820
rect 30984 6808 30990 6860
rect 33520 6857 33548 6888
rect 36998 6876 37004 6888
rect 37056 6876 37062 6928
rect 37185 6919 37243 6925
rect 37185 6885 37197 6919
rect 37231 6916 37243 6919
rect 37366 6916 37372 6928
rect 37231 6888 37372 6916
rect 37231 6885 37243 6888
rect 37185 6879 37243 6885
rect 37366 6876 37372 6888
rect 37424 6876 37430 6928
rect 40052 6888 40356 6916
rect 33505 6851 33563 6857
rect 33505 6817 33517 6851
rect 33551 6817 33563 6851
rect 33505 6811 33563 6817
rect 37550 6808 37556 6860
rect 37608 6848 37614 6860
rect 38289 6851 38347 6857
rect 38289 6848 38301 6851
rect 37608 6820 38301 6848
rect 37608 6808 37614 6820
rect 38289 6817 38301 6820
rect 38335 6817 38347 6851
rect 38289 6811 38347 6817
rect 38470 6808 38476 6860
rect 38528 6848 38534 6860
rect 40052 6848 40080 6888
rect 38528 6820 40080 6848
rect 40328 6848 40356 6888
rect 41874 6876 41880 6928
rect 41932 6916 41938 6928
rect 42337 6919 42395 6925
rect 41932 6888 41977 6916
rect 41932 6876 41938 6888
rect 42337 6885 42349 6919
rect 42383 6885 42395 6919
rect 42337 6879 42395 6885
rect 42812 6888 43116 6916
rect 40865 6851 40923 6857
rect 40865 6848 40877 6851
rect 40328 6820 40877 6848
rect 38528 6808 38534 6820
rect 40865 6817 40877 6820
rect 40911 6817 40923 6851
rect 42352 6848 42380 6879
rect 42812 6857 42840 6888
rect 40865 6811 40923 6817
rect 41616 6820 42380 6848
rect 42797 6851 42855 6857
rect 22097 6783 22155 6789
rect 22097 6780 22109 6783
rect 20416 6684 20484 6712
rect 20548 6752 22109 6780
rect 20416 6681 20428 6684
rect 20370 6675 20428 6681
rect 20548 6656 20576 6752
rect 22097 6749 22109 6752
rect 22143 6749 22155 6783
rect 22278 6780 22284 6792
rect 22239 6752 22284 6780
rect 22097 6743 22155 6749
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 22428 6752 27936 6780
rect 22428 6740 22434 6752
rect 20622 6672 20628 6724
rect 20680 6712 20686 6724
rect 21361 6715 21419 6721
rect 20680 6684 21220 6712
rect 20680 6672 20686 6684
rect 14734 6644 14740 6656
rect 14240 6616 14596 6644
rect 14695 6616 14740 6644
rect 14240 6604 14246 6616
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 16666 6604 16672 6656
rect 16724 6604 16730 6656
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 16942 6644 16948 6656
rect 16807 6616 16948 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 17862 6644 17868 6656
rect 17823 6616 17868 6644
rect 17862 6604 17868 6616
rect 17920 6604 17926 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21192 6653 21220 6684
rect 21361 6681 21373 6715
rect 21407 6712 21419 6715
rect 22462 6712 22468 6724
rect 21407 6684 22468 6712
rect 21407 6681 21419 6684
rect 21361 6675 21419 6681
rect 22462 6672 22468 6684
rect 22520 6672 22526 6724
rect 27908 6712 27936 6752
rect 29546 6740 29552 6792
rect 29604 6780 29610 6792
rect 31018 6780 31024 6792
rect 29604 6752 31024 6780
rect 29604 6740 29610 6752
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 31220 6752 35848 6780
rect 31220 6712 31248 6752
rect 27908 6684 31248 6712
rect 31288 6715 31346 6721
rect 31288 6681 31300 6715
rect 31334 6712 31346 6715
rect 32122 6712 32128 6724
rect 31334 6684 32128 6712
rect 31334 6681 31346 6684
rect 31288 6675 31346 6681
rect 32122 6672 32128 6684
rect 32180 6672 32186 6724
rect 33134 6672 33140 6724
rect 33192 6712 33198 6724
rect 33192 6684 33548 6712
rect 33192 6672 33198 6684
rect 21177 6647 21235 6653
rect 20588 6616 20681 6644
rect 20588 6604 20594 6616
rect 21177 6613 21189 6647
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 21266 6604 21272 6656
rect 21324 6644 21330 6656
rect 21324 6616 21369 6644
rect 21324 6604 21330 6616
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 31386 6644 31392 6656
rect 26292 6616 31392 6644
rect 26292 6604 26298 6616
rect 31386 6604 31392 6616
rect 31444 6604 31450 6656
rect 32398 6644 32404 6656
rect 32359 6616 32404 6644
rect 32398 6604 32404 6616
rect 32456 6644 32462 6656
rect 33226 6644 33232 6656
rect 32456 6616 33232 6644
rect 32456 6604 32462 6616
rect 33226 6604 33232 6616
rect 33284 6604 33290 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 33520 6644 33548 6684
rect 34146 6672 34152 6724
rect 34204 6712 34210 6724
rect 35161 6715 35219 6721
rect 35161 6712 35173 6715
rect 34204 6684 35173 6712
rect 34204 6672 34210 6684
rect 35161 6681 35173 6684
rect 35207 6712 35219 6715
rect 35434 6712 35440 6724
rect 35207 6684 35440 6712
rect 35207 6681 35219 6684
rect 35161 6675 35219 6681
rect 35434 6672 35440 6684
rect 35492 6672 35498 6724
rect 35820 6721 35848 6752
rect 36998 6740 37004 6792
rect 37056 6780 37062 6792
rect 37093 6783 37151 6789
rect 37093 6780 37105 6783
rect 37056 6752 37105 6780
rect 37056 6740 37062 6752
rect 37093 6749 37105 6752
rect 37139 6749 37151 6783
rect 37274 6780 37280 6792
rect 37235 6752 37280 6780
rect 37093 6743 37151 6749
rect 37274 6740 37280 6752
rect 37332 6780 37338 6792
rect 37921 6783 37979 6789
rect 37921 6780 37933 6783
rect 37332 6752 37933 6780
rect 37332 6740 37338 6752
rect 37921 6749 37933 6752
rect 37967 6749 37979 6783
rect 37921 6743 37979 6749
rect 38105 6783 38163 6789
rect 38105 6749 38117 6783
rect 38151 6780 38163 6783
rect 38378 6780 38384 6792
rect 38151 6752 38384 6780
rect 38151 6749 38163 6752
rect 38105 6743 38163 6749
rect 38378 6740 38384 6752
rect 38436 6740 38442 6792
rect 40126 6740 40132 6792
rect 40184 6780 40190 6792
rect 40221 6783 40279 6789
rect 40221 6780 40233 6783
rect 40184 6752 40233 6780
rect 40184 6740 40190 6752
rect 40221 6749 40233 6752
rect 40267 6749 40279 6783
rect 40402 6780 40408 6792
rect 40363 6752 40408 6780
rect 40221 6743 40279 6749
rect 40402 6740 40408 6752
rect 40460 6740 40466 6792
rect 40954 6740 40960 6792
rect 41012 6780 41018 6792
rect 41616 6790 41644 6820
rect 42797 6817 42809 6851
rect 42843 6817 42855 6851
rect 42797 6811 42855 6817
rect 42886 6808 42892 6860
rect 42944 6848 42950 6860
rect 42944 6820 42989 6848
rect 42944 6808 42950 6820
rect 43088 6792 43116 6888
rect 43162 6808 43168 6860
rect 43220 6848 43226 6860
rect 48941 6851 48999 6857
rect 43220 6820 46704 6848
rect 43220 6808 43226 6820
rect 41524 6789 41644 6790
rect 41325 6783 41383 6789
rect 41325 6780 41337 6783
rect 41012 6752 41337 6780
rect 41012 6740 41018 6752
rect 41325 6749 41337 6752
rect 41371 6749 41383 6783
rect 41325 6743 41383 6749
rect 41509 6783 41644 6789
rect 41509 6749 41521 6783
rect 41555 6762 41644 6783
rect 41555 6749 41567 6762
rect 41509 6743 41567 6749
rect 41690 6740 41696 6792
rect 41748 6780 41754 6792
rect 41748 6752 41920 6780
rect 41748 6740 41754 6752
rect 35805 6715 35863 6721
rect 35805 6681 35817 6715
rect 35851 6681 35863 6715
rect 35805 6675 35863 6681
rect 35986 6672 35992 6724
rect 36044 6721 36050 6724
rect 36044 6715 36063 6721
rect 36051 6681 36063 6715
rect 40497 6715 40555 6721
rect 40497 6712 40509 6715
rect 36044 6675 36063 6681
rect 36096 6684 40509 6712
rect 36044 6672 36050 6675
rect 35253 6647 35311 6653
rect 35253 6644 35265 6647
rect 33376 6616 33421 6644
rect 33520 6616 35265 6644
rect 33376 6604 33382 6616
rect 35253 6613 35265 6616
rect 35299 6613 35311 6647
rect 35253 6607 35311 6613
rect 35342 6604 35348 6656
rect 35400 6644 35406 6656
rect 36096 6644 36124 6684
rect 40236 6656 40264 6684
rect 40497 6681 40509 6684
rect 40543 6681 40555 6715
rect 40497 6675 40555 6681
rect 40589 6715 40647 6721
rect 40589 6681 40601 6715
rect 40635 6681 40647 6715
rect 40589 6675 40647 6681
rect 40707 6715 40765 6721
rect 40707 6681 40719 6715
rect 40753 6712 40765 6715
rect 41046 6712 41052 6724
rect 40753 6684 41052 6712
rect 40753 6681 40765 6684
rect 40707 6675 40765 6681
rect 35400 6616 36124 6644
rect 36173 6647 36231 6653
rect 35400 6604 35406 6616
rect 36173 6613 36185 6647
rect 36219 6644 36231 6647
rect 38286 6644 38292 6656
rect 36219 6616 38292 6644
rect 36219 6613 36231 6616
rect 36173 6607 36231 6613
rect 38286 6604 38292 6616
rect 38344 6604 38350 6656
rect 40218 6604 40224 6656
rect 40276 6604 40282 6656
rect 40604 6644 40632 6675
rect 41046 6672 41052 6684
rect 41104 6672 41110 6724
rect 41601 6715 41659 6721
rect 41601 6681 41613 6715
rect 41647 6681 41659 6715
rect 41601 6675 41659 6681
rect 40862 6644 40868 6656
rect 40604 6616 40868 6644
rect 40862 6604 40868 6616
rect 40920 6604 40926 6656
rect 40954 6604 40960 6656
rect 41012 6644 41018 6656
rect 41616 6644 41644 6675
rect 41012 6616 41644 6644
rect 41892 6644 41920 6752
rect 41966 6740 41972 6792
rect 42024 6780 42030 6792
rect 42978 6780 42984 6792
rect 42024 6752 42984 6780
rect 42024 6740 42030 6752
rect 42978 6740 42984 6752
rect 43036 6740 43042 6792
rect 43070 6740 43076 6792
rect 43128 6780 43134 6792
rect 45554 6780 45560 6792
rect 43128 6752 45560 6780
rect 43128 6740 43134 6752
rect 45554 6740 45560 6752
rect 45612 6740 45618 6792
rect 46566 6780 46572 6792
rect 46032 6752 46572 6780
rect 42705 6715 42763 6721
rect 42705 6681 42717 6715
rect 42751 6712 42763 6715
rect 43346 6712 43352 6724
rect 42751 6684 43352 6712
rect 42751 6681 42763 6684
rect 42705 6675 42763 6681
rect 43346 6672 43352 6684
rect 43404 6672 43410 6724
rect 43714 6672 43720 6724
rect 43772 6712 43778 6724
rect 46032 6712 46060 6752
rect 46566 6740 46572 6752
rect 46624 6740 46630 6792
rect 46676 6780 46704 6820
rect 48941 6817 48953 6851
rect 48987 6848 48999 6851
rect 48987 6820 50200 6848
rect 48987 6817 48999 6820
rect 48941 6811 48999 6817
rect 49053 6783 49111 6789
rect 49053 6780 49065 6783
rect 46676 6752 49065 6780
rect 49053 6749 49065 6752
rect 49099 6749 49111 6783
rect 49053 6743 49111 6749
rect 49142 6740 49148 6792
rect 49200 6780 49206 6792
rect 50172 6789 50200 6820
rect 50157 6783 50215 6789
rect 49200 6752 49245 6780
rect 49200 6740 49206 6752
rect 50157 6749 50169 6783
rect 50203 6749 50215 6783
rect 50157 6743 50215 6749
rect 50341 6783 50399 6789
rect 50341 6749 50353 6783
rect 50387 6780 50399 6783
rect 50614 6780 50620 6792
rect 50387 6752 50620 6780
rect 50387 6749 50399 6752
rect 50341 6743 50399 6749
rect 50614 6740 50620 6752
rect 50672 6740 50678 6792
rect 51261 6783 51319 6789
rect 51261 6749 51273 6783
rect 51307 6780 51319 6783
rect 51307 6752 51672 6780
rect 51307 6749 51319 6752
rect 51261 6743 51319 6749
rect 43772 6684 46060 6712
rect 43772 6672 43778 6684
rect 46198 6672 46204 6724
rect 46256 6712 46262 6724
rect 46814 6715 46872 6721
rect 46814 6712 46826 6715
rect 46256 6684 46826 6712
rect 46256 6672 46262 6684
rect 46814 6681 46826 6684
rect 46860 6681 46872 6715
rect 48869 6715 48927 6721
rect 46814 6675 46872 6681
rect 46952 6684 48314 6712
rect 46952 6644 46980 6684
rect 47946 6644 47952 6656
rect 41892 6616 46980 6644
rect 47907 6616 47952 6644
rect 41012 6604 41018 6616
rect 47946 6604 47952 6616
rect 48004 6604 48010 6656
rect 48286 6644 48314 6684
rect 48869 6681 48881 6715
rect 48915 6712 48927 6715
rect 49326 6712 49332 6724
rect 48915 6684 49332 6712
rect 48915 6681 48927 6684
rect 48869 6675 48927 6681
rect 49326 6672 49332 6684
rect 49384 6672 49390 6724
rect 50249 6715 50307 6721
rect 50249 6681 50261 6715
rect 50295 6712 50307 6715
rect 51506 6715 51564 6721
rect 51506 6712 51518 6715
rect 50295 6684 51518 6712
rect 50295 6681 50307 6684
rect 50249 6675 50307 6681
rect 51506 6681 51518 6684
rect 51552 6681 51564 6715
rect 51506 6675 51564 6681
rect 49142 6644 49148 6656
rect 48286 6616 49148 6644
rect 49142 6604 49148 6616
rect 49200 6604 49206 6656
rect 49418 6604 49424 6656
rect 49476 6644 49482 6656
rect 51644 6644 51672 6752
rect 52638 6644 52644 6656
rect 49476 6616 51672 6644
rect 52599 6616 52644 6644
rect 49476 6604 49482 6616
rect 52638 6604 52644 6616
rect 52696 6604 52702 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2774 6440 2780 6452
rect 2735 6412 2780 6440
rect 2774 6400 2780 6412
rect 2832 6400 2838 6452
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 10870 6372 10876 6384
rect 1412 6344 10876 6372
rect 1412 6313 1440 6344
rect 10870 6332 10876 6344
rect 10928 6372 10934 6384
rect 10980 6372 11008 6403
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 17310 6440 17316 6452
rect 15344 6412 17316 6440
rect 15344 6400 15350 6412
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 20073 6443 20131 6449
rect 20073 6409 20085 6443
rect 20119 6440 20131 6443
rect 20162 6440 20168 6452
rect 20119 6412 20168 6440
rect 20119 6409 20131 6412
rect 20073 6403 20131 6409
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 25774 6400 25780 6452
rect 25832 6440 25838 6452
rect 30006 6440 30012 6452
rect 25832 6412 30012 6440
rect 25832 6400 25838 6412
rect 30006 6400 30012 6412
rect 30064 6400 30070 6452
rect 30291 6443 30349 6449
rect 30291 6440 30303 6443
rect 30116 6412 30303 6440
rect 10928 6344 11008 6372
rect 10928 6332 10934 6344
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 20809 6375 20867 6381
rect 20809 6372 20821 6375
rect 20036 6344 20821 6372
rect 20036 6332 20042 6344
rect 20809 6341 20821 6344
rect 20855 6341 20867 6375
rect 24394 6372 24400 6384
rect 20809 6335 20867 6341
rect 22757 6344 24400 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2958 6304 2964 6316
rect 2363 6276 2964 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 5166 6304 5172 6316
rect 3191 6276 5172 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 9858 6313 9864 6316
rect 9852 6267 9864 6313
rect 9916 6304 9922 6316
rect 9916 6276 9952 6304
rect 9858 6264 9864 6267
rect 9916 6264 9922 6276
rect 10594 6264 10600 6316
rect 10652 6304 10658 6316
rect 13262 6304 13268 6316
rect 10652 6276 13268 6304
rect 10652 6264 10658 6276
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 16264 6276 17417 6304
rect 16264 6264 16270 6276
rect 17405 6273 17417 6276
rect 17451 6304 17463 6307
rect 19426 6304 19432 6316
rect 17451 6276 19432 6304
rect 17451 6273 17463 6276
rect 17405 6267 17463 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 20530 6304 20536 6316
rect 19751 6276 20536 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 21450 6264 21456 6316
rect 21508 6304 21514 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21508 6276 22017 6304
rect 21508 6264 21514 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 22757 6304 22785 6344
rect 24394 6332 24400 6344
rect 24452 6332 24458 6384
rect 29472 6344 29776 6372
rect 22235 6276 22785 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 22830 6264 22836 6316
rect 22888 6304 22894 6316
rect 25866 6304 25872 6316
rect 22888 6276 25872 6304
rect 22888 6264 22894 6276
rect 25866 6264 25872 6276
rect 25924 6264 25930 6316
rect 26050 6304 26056 6316
rect 26011 6276 26056 6304
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 26234 6304 26240 6316
rect 26195 6276 26240 6304
rect 26234 6264 26240 6276
rect 26292 6264 26298 6316
rect 26786 6264 26792 6316
rect 26844 6304 26850 6316
rect 29086 6304 29092 6316
rect 26844 6276 29092 6304
rect 26844 6264 26850 6276
rect 29086 6264 29092 6276
rect 29144 6264 29150 6316
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 2648 6208 3341 6236
rect 2648 6196 2654 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 3329 6199 3387 6205
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 11940 6208 17141 6236
rect 11940 6196 11946 6208
rect 17129 6205 17141 6208
rect 17175 6236 17187 6239
rect 20806 6236 20812 6248
rect 17175 6208 20812 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 22094 6196 22100 6248
rect 22152 6236 22158 6248
rect 22278 6236 22284 6248
rect 22152 6208 22197 6236
rect 22239 6208 22284 6236
rect 22152 6196 22158 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22462 6196 22468 6248
rect 22520 6236 22526 6248
rect 26252 6236 26280 6264
rect 29472 6236 29500 6344
rect 29748 6316 29776 6344
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6273 29607 6307
rect 29730 6304 29736 6316
rect 29691 6276 29736 6304
rect 29549 6267 29607 6273
rect 22520 6208 26280 6236
rect 28966 6208 29500 6236
rect 29564 6236 29592 6267
rect 29730 6264 29736 6276
rect 29788 6264 29794 6316
rect 30116 6304 30144 6412
rect 30291 6409 30303 6412
rect 30337 6409 30349 6443
rect 30291 6403 30349 6409
rect 30377 6443 30435 6449
rect 30377 6409 30389 6443
rect 30423 6440 30435 6443
rect 31110 6440 31116 6452
rect 30423 6412 31116 6440
rect 30423 6409 30435 6412
rect 30377 6403 30435 6409
rect 31110 6400 31116 6412
rect 31168 6400 31174 6452
rect 33318 6440 33324 6452
rect 31220 6412 33324 6440
rect 30193 6375 30251 6381
rect 30193 6341 30205 6375
rect 30239 6372 30251 6375
rect 30650 6372 30656 6384
rect 30239 6344 30656 6372
rect 30239 6341 30251 6344
rect 30193 6335 30251 6341
rect 30650 6332 30656 6344
rect 30708 6332 30714 6384
rect 30926 6332 30932 6384
rect 30984 6372 30990 6384
rect 31220 6372 31248 6412
rect 33318 6400 33324 6412
rect 33376 6400 33382 6452
rect 36078 6440 36084 6452
rect 33428 6412 36084 6440
rect 30984 6344 31248 6372
rect 30984 6332 30990 6344
rect 32214 6332 32220 6384
rect 32272 6372 32278 6384
rect 33428 6372 33456 6412
rect 36078 6400 36084 6412
rect 36136 6400 36142 6452
rect 36262 6400 36268 6452
rect 36320 6440 36326 6452
rect 36320 6412 38792 6440
rect 36320 6400 36326 6412
rect 37734 6372 37740 6384
rect 32272 6344 33456 6372
rect 35084 6344 37740 6372
rect 32272 6332 32278 6344
rect 30466 6304 30472 6316
rect 29840 6276 30144 6304
rect 30427 6276 30472 6304
rect 29840 6236 29868 6276
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 31018 6264 31024 6316
rect 31076 6304 31082 6316
rect 33410 6304 33416 6316
rect 31076 6276 33416 6304
rect 31076 6264 31082 6276
rect 33410 6264 33416 6276
rect 33468 6264 33474 6316
rect 34146 6304 34152 6316
rect 34107 6276 34152 6304
rect 34146 6264 34152 6276
rect 34204 6264 34210 6316
rect 34238 6264 34244 6316
rect 34296 6304 34302 6316
rect 35084 6313 35112 6344
rect 37734 6332 37740 6344
rect 37792 6332 37798 6384
rect 38473 6375 38531 6381
rect 38473 6341 38485 6375
rect 38519 6372 38531 6375
rect 38562 6372 38568 6384
rect 38519 6344 38568 6372
rect 38519 6341 38531 6344
rect 38473 6335 38531 6341
rect 38562 6332 38568 6344
rect 38620 6332 38626 6384
rect 38764 6372 38792 6412
rect 40402 6400 40408 6452
rect 40460 6440 40466 6452
rect 42797 6443 42855 6449
rect 42797 6440 42809 6443
rect 40460 6412 42809 6440
rect 40460 6400 40466 6412
rect 42797 6409 42809 6412
rect 42843 6409 42855 6443
rect 46934 6440 46940 6452
rect 46895 6412 46940 6440
rect 42797 6403 42855 6409
rect 46934 6400 46940 6412
rect 46992 6400 46998 6452
rect 47026 6400 47032 6452
rect 47084 6440 47090 6452
rect 48866 6440 48872 6452
rect 47084 6412 48872 6440
rect 47084 6400 47090 6412
rect 48866 6400 48872 6412
rect 48924 6400 48930 6452
rect 38764 6344 39528 6372
rect 35069 6307 35127 6313
rect 35069 6304 35081 6307
rect 34296 6276 35081 6304
rect 34296 6264 34302 6276
rect 35069 6273 35081 6276
rect 35115 6273 35127 6307
rect 35069 6267 35127 6273
rect 35253 6307 35311 6313
rect 35253 6273 35265 6307
rect 35299 6304 35311 6307
rect 35342 6304 35348 6316
rect 35299 6276 35348 6304
rect 35299 6273 35311 6276
rect 35253 6267 35311 6273
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 36265 6307 36323 6313
rect 36265 6273 36277 6307
rect 36311 6304 36323 6307
rect 36354 6304 36360 6316
rect 36311 6276 36360 6304
rect 36311 6273 36323 6276
rect 36265 6267 36323 6273
rect 34790 6236 34796 6248
rect 29564 6208 29868 6236
rect 31726 6208 34796 6236
rect 22520 6196 22526 6208
rect 2133 6171 2191 6177
rect 2133 6137 2145 6171
rect 2179 6168 2191 6171
rect 8294 6168 8300 6180
rect 2179 6140 8300 6168
rect 2179 6137 2191 6140
rect 2133 6131 2191 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 19306 6140 20668 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 14274 6100 14280 6112
rect 8904 6072 14280 6100
rect 8904 6060 8910 6072
rect 14274 6060 14280 6072
rect 14332 6100 14338 6112
rect 19306 6100 19334 6140
rect 14332 6072 19334 6100
rect 14332 6060 14338 6072
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 20036 6072 20085 6100
rect 20036 6060 20042 6072
rect 20073 6069 20085 6072
rect 20119 6069 20131 6103
rect 20254 6100 20260 6112
rect 20215 6072 20260 6100
rect 20073 6063 20131 6069
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 20640 6100 20668 6140
rect 20714 6128 20720 6180
rect 20772 6168 20778 6180
rect 21085 6171 21143 6177
rect 21085 6168 21097 6171
rect 20772 6140 21097 6168
rect 20772 6128 20778 6140
rect 21085 6137 21097 6140
rect 21131 6168 21143 6171
rect 21131 6140 22094 6168
rect 21131 6137 21143 6140
rect 21085 6131 21143 6137
rect 21634 6100 21640 6112
rect 20640 6072 21640 6100
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 22066 6100 22094 6140
rect 22186 6128 22192 6180
rect 22244 6168 22250 6180
rect 28966 6168 28994 6208
rect 31726 6168 31754 6208
rect 34790 6196 34796 6208
rect 34848 6196 34854 6248
rect 35986 6196 35992 6248
rect 36044 6236 36050 6248
rect 36280 6236 36308 6267
rect 36354 6264 36360 6276
rect 36412 6264 36418 6316
rect 36906 6264 36912 6316
rect 36964 6304 36970 6316
rect 38764 6313 38792 6344
rect 38657 6307 38715 6313
rect 38657 6304 38669 6307
rect 36964 6276 38669 6304
rect 36964 6264 36970 6276
rect 38657 6273 38669 6276
rect 38703 6273 38715 6307
rect 38657 6267 38715 6273
rect 38749 6307 38807 6313
rect 38749 6273 38761 6307
rect 38795 6273 38807 6307
rect 38749 6267 38807 6273
rect 39209 6307 39267 6313
rect 39209 6273 39221 6307
rect 39255 6273 39267 6307
rect 39390 6304 39396 6316
rect 39351 6276 39396 6304
rect 39209 6267 39267 6273
rect 39224 6236 39252 6267
rect 39390 6264 39396 6276
rect 39448 6264 39454 6316
rect 39500 6304 39528 6344
rect 40126 6332 40132 6384
rect 40184 6372 40190 6384
rect 44238 6375 44296 6381
rect 44238 6372 44250 6375
rect 40184 6344 42288 6372
rect 40184 6332 40190 6344
rect 41141 6307 41199 6313
rect 39500 6276 41092 6304
rect 36044 6208 36308 6236
rect 38488 6208 39252 6236
rect 36044 6196 36050 6208
rect 22244 6140 28994 6168
rect 29472 6140 31754 6168
rect 22244 6128 22250 6140
rect 22462 6100 22468 6112
rect 22066 6072 22468 6100
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 25590 6060 25596 6112
rect 25648 6100 25654 6112
rect 26053 6103 26111 6109
rect 26053 6100 26065 6103
rect 25648 6072 26065 6100
rect 25648 6060 25654 6072
rect 26053 6069 26065 6072
rect 26099 6069 26111 6103
rect 26053 6063 26111 6069
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 29472 6100 29500 6140
rect 33686 6128 33692 6180
rect 33744 6168 33750 6180
rect 38488 6177 38516 6208
rect 40862 6196 40868 6248
rect 40920 6236 40926 6248
rect 40957 6239 41015 6245
rect 40957 6236 40969 6239
rect 40920 6208 40969 6236
rect 40920 6196 40926 6208
rect 40957 6205 40969 6208
rect 41003 6205 41015 6239
rect 41064 6236 41092 6276
rect 41141 6273 41153 6307
rect 41187 6304 41199 6307
rect 41874 6304 41880 6316
rect 41187 6276 41880 6304
rect 41187 6273 41199 6276
rect 41141 6267 41199 6273
rect 41874 6264 41880 6276
rect 41932 6264 41938 6316
rect 42260 6304 42288 6344
rect 42996 6344 44250 6372
rect 42996 6304 43024 6344
rect 44238 6341 44250 6344
rect 44284 6341 44296 6375
rect 44238 6335 44296 6341
rect 47581 6375 47639 6381
rect 47581 6341 47593 6375
rect 47627 6372 47639 6375
rect 49022 6375 49080 6381
rect 49022 6372 49034 6375
rect 47627 6344 49034 6372
rect 47627 6341 47639 6344
rect 47581 6335 47639 6341
rect 49022 6341 49034 6344
rect 49068 6341 49080 6375
rect 49022 6335 49080 6341
rect 42260 6276 43024 6304
rect 43070 6264 43076 6316
rect 43128 6304 43134 6316
rect 43165 6307 43223 6313
rect 43165 6304 43177 6307
rect 43128 6276 43177 6304
rect 43128 6264 43134 6276
rect 43165 6273 43177 6276
rect 43211 6273 43223 6307
rect 43165 6267 43223 6273
rect 43530 6264 43536 6316
rect 43588 6304 43594 6316
rect 46385 6307 46443 6313
rect 46385 6304 46397 6307
rect 43588 6276 46397 6304
rect 43588 6264 43594 6276
rect 46385 6273 46397 6276
rect 46431 6273 46443 6307
rect 46566 6304 46572 6316
rect 46527 6276 46572 6304
rect 46385 6267 46443 6273
rect 46566 6264 46572 6276
rect 46624 6264 46630 6316
rect 46658 6264 46664 6316
rect 46716 6304 46722 6316
rect 46799 6307 46857 6313
rect 46716 6276 46761 6304
rect 46716 6264 46722 6276
rect 46799 6273 46811 6307
rect 46845 6304 46857 6307
rect 47118 6304 47124 6316
rect 46845 6276 47124 6304
rect 46845 6273 46857 6276
rect 46799 6267 46857 6273
rect 47118 6264 47124 6276
rect 47176 6264 47182 6316
rect 47302 6264 47308 6316
rect 47360 6304 47366 6316
rect 47765 6307 47823 6313
rect 47765 6304 47777 6307
rect 47360 6276 47777 6304
rect 47360 6264 47366 6276
rect 47765 6273 47777 6276
rect 47811 6273 47823 6307
rect 47765 6267 47823 6273
rect 41598 6236 41604 6248
rect 41064 6208 41604 6236
rect 40957 6199 41015 6205
rect 41598 6196 41604 6208
rect 41656 6196 41662 6248
rect 43254 6236 43260 6248
rect 43215 6208 43260 6236
rect 43254 6196 43260 6208
rect 43312 6196 43318 6248
rect 43349 6239 43407 6245
rect 43349 6205 43361 6239
rect 43395 6205 43407 6239
rect 43349 6199 43407 6205
rect 38473 6171 38531 6177
rect 33744 6140 35204 6168
rect 33744 6128 33750 6140
rect 26200 6072 29500 6100
rect 29549 6103 29607 6109
rect 26200 6060 26206 6072
rect 29549 6069 29561 6103
rect 29595 6100 29607 6103
rect 29638 6100 29644 6112
rect 29595 6072 29644 6100
rect 29595 6069 29607 6072
rect 29549 6063 29607 6069
rect 29638 6060 29644 6072
rect 29696 6060 29702 6112
rect 34422 6060 34428 6112
rect 34480 6100 34486 6112
rect 34480 6072 34525 6100
rect 34480 6060 34486 6072
rect 34698 6060 34704 6112
rect 34756 6100 34762 6112
rect 35069 6103 35127 6109
rect 35069 6100 35081 6103
rect 34756 6072 35081 6100
rect 34756 6060 34762 6072
rect 35069 6069 35081 6072
rect 35115 6069 35127 6103
rect 35176 6100 35204 6140
rect 38473 6137 38485 6171
rect 38519 6137 38531 6171
rect 38473 6131 38531 6137
rect 38562 6128 38568 6180
rect 38620 6168 38626 6180
rect 39390 6168 39396 6180
rect 38620 6140 39396 6168
rect 38620 6128 38626 6140
rect 39390 6128 39396 6140
rect 39448 6128 39454 6180
rect 42702 6128 42708 6180
rect 42760 6168 42766 6180
rect 43364 6168 43392 6199
rect 43714 6196 43720 6248
rect 43772 6236 43778 6248
rect 43993 6239 44051 6245
rect 43993 6236 44005 6239
rect 43772 6208 44005 6236
rect 43772 6196 43778 6208
rect 43993 6205 44005 6208
rect 44039 6205 44051 6239
rect 48038 6236 48044 6248
rect 47999 6208 48044 6236
rect 43993 6199 44051 6205
rect 48038 6196 48044 6208
rect 48096 6196 48102 6248
rect 48777 6239 48835 6245
rect 48777 6205 48789 6239
rect 48823 6205 48835 6239
rect 48777 6199 48835 6205
rect 47949 6171 48007 6177
rect 47949 6168 47961 6171
rect 42760 6140 43392 6168
rect 44928 6140 47961 6168
rect 42760 6128 42766 6140
rect 36357 6103 36415 6109
rect 36357 6100 36369 6103
rect 35176 6072 36369 6100
rect 35069 6063 35127 6069
rect 36357 6069 36369 6072
rect 36403 6100 36415 6103
rect 36722 6100 36728 6112
rect 36403 6072 36728 6100
rect 36403 6069 36415 6072
rect 36357 6063 36415 6069
rect 36722 6060 36728 6072
rect 36780 6060 36786 6112
rect 39206 6100 39212 6112
rect 39167 6072 39212 6100
rect 39206 6060 39212 6072
rect 39264 6060 39270 6112
rect 41325 6103 41383 6109
rect 41325 6069 41337 6103
rect 41371 6100 41383 6103
rect 41506 6100 41512 6112
rect 41371 6072 41512 6100
rect 41371 6069 41383 6072
rect 41325 6063 41383 6069
rect 41506 6060 41512 6072
rect 41564 6060 41570 6112
rect 41690 6060 41696 6112
rect 41748 6100 41754 6112
rect 44928 6100 44956 6140
rect 47949 6137 47961 6140
rect 47995 6137 48007 6171
rect 47949 6131 48007 6137
rect 41748 6072 44956 6100
rect 45373 6103 45431 6109
rect 41748 6060 41754 6072
rect 45373 6069 45385 6103
rect 45419 6100 45431 6103
rect 45554 6100 45560 6112
rect 45419 6072 45560 6100
rect 45419 6069 45431 6072
rect 45373 6063 45431 6069
rect 45554 6060 45560 6072
rect 45612 6100 45618 6112
rect 46750 6100 46756 6112
rect 45612 6072 46756 6100
rect 45612 6060 45618 6072
rect 46750 6060 46756 6072
rect 46808 6060 46814 6112
rect 46842 6060 46848 6112
rect 46900 6100 46906 6112
rect 48590 6100 48596 6112
rect 46900 6072 48596 6100
rect 46900 6060 46906 6072
rect 48590 6060 48596 6072
rect 48648 6100 48654 6112
rect 48792 6100 48820 6199
rect 49418 6100 49424 6112
rect 48648 6072 49424 6100
rect 48648 6060 48654 6072
rect 49418 6060 49424 6072
rect 49476 6060 49482 6112
rect 50154 6100 50160 6112
rect 50115 6072 50160 6100
rect 50154 6060 50160 6072
rect 50212 6060 50218 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 7834 5896 7840 5908
rect 7795 5868 7840 5896
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9916 5868 9965 5896
rect 9916 5856 9922 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 19978 5896 19984 5908
rect 19939 5868 19984 5896
rect 9953 5859 10011 5865
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 22186 5896 22192 5908
rect 20680 5868 22192 5896
rect 20680 5856 20686 5868
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 41874 5896 41880 5908
rect 22296 5868 41880 5896
rect 2608 5800 4384 5828
rect 2608 5772 2636 5800
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2648 5732 2693 5760
rect 2648 5720 2654 5732
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4356 5769 4384 5800
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 13078 5828 13084 5840
rect 12492 5800 13084 5828
rect 12492 5788 12498 5800
rect 13078 5788 13084 5800
rect 13136 5828 13142 5840
rect 19886 5828 19892 5840
rect 13136 5800 19892 5828
rect 13136 5788 13142 5800
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 21450 5828 21456 5840
rect 21411 5800 21456 5828
rect 21450 5788 21456 5800
rect 21508 5788 21514 5840
rect 22005 5831 22063 5837
rect 22005 5797 22017 5831
rect 22051 5828 22063 5831
rect 22094 5828 22100 5840
rect 22051 5800 22100 5828
rect 22051 5797 22063 5800
rect 22005 5791 22063 5797
rect 22094 5788 22100 5800
rect 22152 5788 22158 5840
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 3660 5732 4261 5760
rect 3660 5720 3666 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 20622 5760 20628 5772
rect 11112 5732 20628 5760
rect 11112 5720 11118 5732
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 21726 5720 21732 5772
rect 21784 5760 21790 5772
rect 22296 5760 22324 5868
rect 41874 5856 41880 5868
rect 41932 5856 41938 5908
rect 47302 5896 47308 5908
rect 41984 5868 47308 5896
rect 27614 5828 27620 5840
rect 27575 5800 27620 5828
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 30926 5828 30932 5840
rect 30887 5800 30932 5828
rect 30926 5788 30932 5800
rect 30984 5788 30990 5840
rect 31956 5800 32352 5828
rect 21784 5732 22324 5760
rect 21784 5720 21790 5732
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 24118 5760 24124 5772
rect 23532 5732 24124 5760
rect 23532 5720 23538 5732
rect 24118 5720 24124 5732
rect 24176 5760 24182 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 24176 5732 24409 5760
rect 24176 5720 24182 5732
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 3142 5692 3148 5704
rect 1627 5664 3148 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 6086 5652 6092 5704
rect 6144 5692 6150 5704
rect 6457 5695 6515 5701
rect 6457 5692 6469 5695
rect 6144 5664 6469 5692
rect 6144 5652 6150 5664
rect 6457 5661 6469 5664
rect 6503 5661 6515 5695
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 6457 5655 6515 5661
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10376 5664 10425 5692
rect 10376 5652 10382 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13872 5664 14289 5692
rect 13872 5652 13878 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 14277 5655 14335 5661
rect 4246 5624 4252 5636
rect 2056 5596 4252 5624
rect 2056 5565 2084 5596
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 6724 5627 6782 5633
rect 6724 5593 6736 5627
rect 6770 5624 6782 5627
rect 7926 5624 7932 5636
rect 6770 5596 7932 5624
rect 6770 5593 6782 5596
rect 6724 5587 6782 5593
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 12894 5624 12900 5636
rect 9548 5596 12900 5624
rect 9548 5584 9554 5596
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 2041 5559 2099 5565
rect 2041 5525 2053 5559
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 3326 5556 3332 5568
rect 2455 5528 3332 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 3602 5516 3608 5568
rect 3660 5556 3666 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3660 5528 3801 5556
rect 3660 5516 3666 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5556 4215 5559
rect 5166 5556 5172 5568
rect 4203 5528 5172 5556
rect 4203 5525 4215 5528
rect 4157 5519 4215 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 10321 5559 10379 5565
rect 10321 5556 10333 5559
rect 7248 5528 10333 5556
rect 7248 5516 7254 5528
rect 10321 5525 10333 5528
rect 10367 5525 10379 5559
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 10321 5519 10379 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14292 5556 14320 5655
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 16390 5692 16396 5704
rect 14599 5664 16396 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 16390 5652 16396 5664
rect 16448 5652 16454 5704
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20162 5692 20168 5704
rect 20036 5664 20168 5692
rect 20036 5652 20042 5664
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 21085 5695 21143 5701
rect 21085 5692 21097 5695
rect 20487 5664 21097 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 21085 5661 21097 5664
rect 21131 5692 21143 5695
rect 21910 5692 21916 5704
rect 21131 5664 21916 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22097 5695 22155 5701
rect 22097 5661 22109 5695
rect 22143 5661 22155 5695
rect 24412 5692 24440 5723
rect 29086 5720 29092 5772
rect 29144 5760 29150 5772
rect 29546 5760 29552 5772
rect 29144 5732 29552 5760
rect 29144 5720 29150 5732
rect 29546 5720 29552 5732
rect 29604 5720 29610 5772
rect 26237 5695 26295 5701
rect 26237 5692 26249 5695
rect 24412 5664 26249 5692
rect 22097 5655 22155 5661
rect 26237 5661 26249 5664
rect 26283 5692 26295 5695
rect 26786 5692 26792 5704
rect 26283 5664 26792 5692
rect 26283 5661 26295 5664
rect 26237 5655 26295 5661
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 20349 5627 20407 5633
rect 20349 5624 20361 5627
rect 19484 5596 20361 5624
rect 19484 5584 19490 5596
rect 20349 5593 20361 5596
rect 20395 5624 20407 5627
rect 21269 5627 21327 5633
rect 21269 5624 21281 5627
rect 20395 5596 21281 5624
rect 20395 5593 20407 5596
rect 20349 5587 20407 5593
rect 21269 5593 21281 5596
rect 21315 5593 21327 5627
rect 21269 5587 21327 5593
rect 21174 5556 21180 5568
rect 14292 5528 21180 5556
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 21284 5556 21312 5587
rect 22112 5556 22140 5655
rect 26786 5652 26792 5664
rect 26844 5652 26850 5704
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 29805 5695 29863 5701
rect 29805 5692 29817 5695
rect 29696 5664 29817 5692
rect 29696 5652 29702 5664
rect 29805 5661 29817 5664
rect 29851 5661 29863 5695
rect 29805 5655 29863 5661
rect 24664 5627 24722 5633
rect 24664 5593 24676 5627
rect 24710 5624 24722 5627
rect 24854 5624 24860 5636
rect 24710 5596 24860 5624
rect 24710 5593 24722 5596
rect 24664 5587 24722 5593
rect 24854 5584 24860 5596
rect 24912 5584 24918 5636
rect 26326 5584 26332 5636
rect 26384 5624 26390 5636
rect 26482 5627 26540 5633
rect 26482 5624 26494 5627
rect 26384 5596 26494 5624
rect 26384 5584 26390 5596
rect 26482 5593 26494 5596
rect 26528 5593 26540 5627
rect 26482 5587 26540 5593
rect 26970 5584 26976 5636
rect 27028 5624 27034 5636
rect 31956 5624 31984 5800
rect 32214 5720 32220 5772
rect 32272 5720 32278 5772
rect 32324 5760 32352 5800
rect 33042 5788 33048 5840
rect 33100 5828 33106 5840
rect 34698 5828 34704 5840
rect 33100 5800 34704 5828
rect 33100 5788 33106 5800
rect 34698 5788 34704 5800
rect 34756 5788 34762 5840
rect 35526 5788 35532 5840
rect 35584 5828 35590 5840
rect 35713 5831 35771 5837
rect 35713 5828 35725 5831
rect 35584 5800 35725 5828
rect 35584 5788 35590 5800
rect 35713 5797 35725 5800
rect 35759 5797 35771 5831
rect 41984 5828 42012 5868
rect 47302 5856 47308 5868
rect 47360 5856 47366 5908
rect 47486 5856 47492 5908
rect 47544 5896 47550 5908
rect 50614 5896 50620 5908
rect 47544 5868 50620 5896
rect 47544 5856 47550 5868
rect 43346 5828 43352 5840
rect 35713 5791 35771 5797
rect 35820 5800 42012 5828
rect 43307 5800 43352 5828
rect 35820 5760 35848 5800
rect 43346 5788 43352 5800
rect 43404 5788 43410 5840
rect 47026 5828 47032 5840
rect 44928 5800 47032 5828
rect 32324 5732 35848 5760
rect 35912 5732 42104 5760
rect 32033 5695 32091 5701
rect 32033 5661 32045 5695
rect 32079 5661 32091 5695
rect 32033 5655 32091 5661
rect 32125 5695 32183 5701
rect 32125 5661 32137 5695
rect 32171 5692 32183 5695
rect 32232 5692 32260 5720
rect 34698 5692 34704 5704
rect 32171 5664 32260 5692
rect 34659 5664 34704 5692
rect 32171 5661 32183 5664
rect 32125 5655 32183 5661
rect 27028 5596 31984 5624
rect 32048 5624 32076 5655
rect 34698 5652 34704 5664
rect 34756 5652 34762 5704
rect 34885 5695 34943 5701
rect 34885 5661 34897 5695
rect 34931 5661 34943 5695
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 34885 5655 34943 5661
rect 34992 5664 35725 5692
rect 33134 5624 33140 5636
rect 32048 5596 33140 5624
rect 27028 5584 27034 5596
rect 33134 5584 33140 5596
rect 33192 5624 33198 5636
rect 34900 5624 34928 5655
rect 33192 5596 34928 5624
rect 33192 5584 33198 5596
rect 21284 5528 22140 5556
rect 25777 5559 25835 5565
rect 25777 5525 25789 5559
rect 25823 5556 25835 5559
rect 25866 5556 25872 5568
rect 25823 5528 25872 5556
rect 25823 5525 25835 5528
rect 25777 5519 25835 5525
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 26050 5516 26056 5568
rect 26108 5556 26114 5568
rect 32033 5559 32091 5565
rect 32033 5556 32045 5559
rect 26108 5528 32045 5556
rect 26108 5516 26114 5528
rect 32033 5525 32045 5528
rect 32079 5525 32091 5559
rect 32033 5519 32091 5525
rect 32490 5516 32496 5568
rect 32548 5556 32554 5568
rect 34992 5556 35020 5664
rect 35713 5661 35725 5664
rect 35759 5692 35771 5695
rect 35912 5692 35940 5732
rect 35759 5664 35940 5692
rect 35989 5695 36047 5701
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 35989 5661 36001 5695
rect 36035 5692 36047 5695
rect 36354 5692 36360 5704
rect 36035 5664 36360 5692
rect 36035 5661 36047 5664
rect 35989 5655 36047 5661
rect 36354 5652 36360 5664
rect 36412 5652 36418 5704
rect 38194 5652 38200 5704
rect 38252 5692 38258 5704
rect 41230 5692 41236 5704
rect 38252 5664 41236 5692
rect 38252 5652 38258 5664
rect 41230 5652 41236 5664
rect 41288 5652 41294 5704
rect 41506 5692 41512 5704
rect 41467 5664 41512 5692
rect 41506 5652 41512 5664
rect 41564 5652 41570 5704
rect 41966 5692 41972 5704
rect 41927 5664 41972 5692
rect 41966 5652 41972 5664
rect 42024 5652 42030 5704
rect 42076 5692 42104 5732
rect 43254 5720 43260 5772
rect 43312 5760 43318 5772
rect 44928 5760 44956 5800
rect 47026 5788 47032 5800
rect 47084 5788 47090 5840
rect 47397 5831 47455 5837
rect 47397 5797 47409 5831
rect 47443 5828 47455 5831
rect 48038 5828 48044 5840
rect 47443 5800 48044 5828
rect 47443 5797 47455 5800
rect 47397 5791 47455 5797
rect 48038 5788 48044 5800
rect 48096 5788 48102 5840
rect 48777 5831 48835 5837
rect 48777 5797 48789 5831
rect 48823 5797 48835 5831
rect 48777 5791 48835 5797
rect 46566 5760 46572 5772
rect 43312 5732 44956 5760
rect 45020 5732 46572 5760
rect 43312 5720 43318 5732
rect 45020 5692 45048 5732
rect 46566 5720 46572 5732
rect 46624 5760 46630 5772
rect 46624 5732 46980 5760
rect 46624 5720 46630 5732
rect 42076 5664 45048 5692
rect 45094 5652 45100 5704
rect 45152 5692 45158 5704
rect 45152 5664 45197 5692
rect 45152 5652 45158 5664
rect 46658 5652 46664 5704
rect 46716 5692 46722 5704
rect 46845 5695 46903 5701
rect 46845 5692 46857 5695
rect 46716 5664 46857 5692
rect 46716 5652 46722 5664
rect 46845 5661 46857 5664
rect 46891 5661 46903 5695
rect 46845 5655 46903 5661
rect 35158 5584 35164 5636
rect 35216 5624 35222 5636
rect 35894 5624 35900 5636
rect 35216 5596 35572 5624
rect 35855 5596 35900 5624
rect 35216 5584 35222 5596
rect 32548 5528 35020 5556
rect 35069 5559 35127 5565
rect 32548 5516 32554 5528
rect 35069 5525 35081 5559
rect 35115 5556 35127 5559
rect 35434 5556 35440 5568
rect 35115 5528 35440 5556
rect 35115 5525 35127 5528
rect 35069 5519 35127 5525
rect 35434 5516 35440 5528
rect 35492 5516 35498 5568
rect 35544 5556 35572 5596
rect 35894 5584 35900 5596
rect 35952 5584 35958 5636
rect 36722 5584 36728 5636
rect 36780 5624 36786 5636
rect 40218 5624 40224 5636
rect 36780 5596 40224 5624
rect 36780 5584 36786 5596
rect 40218 5584 40224 5596
rect 40276 5584 40282 5636
rect 40313 5627 40371 5633
rect 40313 5593 40325 5627
rect 40359 5624 40371 5627
rect 40402 5624 40408 5636
rect 40359 5596 40408 5624
rect 40359 5593 40371 5596
rect 40313 5587 40371 5593
rect 40402 5584 40408 5596
rect 40460 5584 40466 5636
rect 40497 5627 40555 5633
rect 40497 5593 40509 5627
rect 40543 5624 40555 5627
rect 40862 5624 40868 5636
rect 40543 5596 40868 5624
rect 40543 5593 40555 5596
rect 40497 5587 40555 5593
rect 40862 5584 40868 5596
rect 40920 5584 40926 5636
rect 42214 5627 42272 5633
rect 42214 5624 42226 5627
rect 41340 5596 42226 5624
rect 40954 5556 40960 5568
rect 35544 5528 40960 5556
rect 40954 5516 40960 5528
rect 41012 5516 41018 5568
rect 41340 5565 41368 5596
rect 42214 5593 42226 5596
rect 42260 5593 42272 5627
rect 45646 5624 45652 5636
rect 42214 5587 42272 5593
rect 43732 5596 45652 5624
rect 43732 5568 43760 5596
rect 45646 5584 45652 5596
rect 45704 5584 45710 5636
rect 41325 5559 41383 5565
rect 41325 5525 41337 5559
rect 41371 5525 41383 5559
rect 41325 5519 41383 5525
rect 41966 5516 41972 5568
rect 42024 5556 42030 5568
rect 43714 5556 43720 5568
rect 42024 5528 43720 5556
rect 42024 5516 42030 5528
rect 43714 5516 43720 5528
rect 43772 5516 43778 5568
rect 45278 5556 45284 5568
rect 45239 5528 45284 5556
rect 45278 5516 45284 5528
rect 45336 5516 45342 5568
rect 46860 5556 46888 5655
rect 46952 5624 46980 5732
rect 47118 5720 47124 5772
rect 47176 5720 47182 5772
rect 48792 5760 48820 5791
rect 48792 5732 50200 5760
rect 47136 5692 47164 5720
rect 47237 5695 47295 5701
rect 47237 5692 47249 5695
rect 47136 5664 47249 5692
rect 47237 5661 47249 5664
rect 47283 5661 47295 5695
rect 47237 5655 47295 5661
rect 47394 5652 47400 5704
rect 47452 5692 47458 5704
rect 48961 5695 49019 5701
rect 48961 5692 48973 5695
rect 47452 5664 48973 5692
rect 47452 5652 47458 5664
rect 48961 5661 48973 5664
rect 49007 5661 49019 5695
rect 48961 5655 49019 5661
rect 49053 5695 49111 5701
rect 49053 5661 49065 5695
rect 49099 5692 49111 5695
rect 49142 5692 49148 5704
rect 49099 5664 49148 5692
rect 49099 5661 49111 5664
rect 49053 5655 49111 5661
rect 49142 5652 49148 5664
rect 49200 5652 49206 5704
rect 50172 5701 50200 5732
rect 50157 5695 50215 5701
rect 50157 5661 50169 5695
rect 50203 5661 50215 5695
rect 50264 5692 50292 5868
rect 50614 5856 50620 5868
rect 50672 5856 50678 5908
rect 50341 5695 50399 5701
rect 50341 5692 50353 5695
rect 50264 5664 50353 5692
rect 50157 5655 50215 5661
rect 50341 5661 50353 5664
rect 50387 5661 50399 5695
rect 50341 5655 50399 5661
rect 47026 5624 47032 5636
rect 46939 5596 47032 5624
rect 47026 5584 47032 5596
rect 47084 5584 47090 5636
rect 47121 5627 47179 5633
rect 47121 5593 47133 5627
rect 47167 5624 47179 5627
rect 48774 5624 48780 5636
rect 47167 5596 48636 5624
rect 48735 5596 48780 5624
rect 47167 5593 47179 5596
rect 47121 5587 47179 5593
rect 47946 5556 47952 5568
rect 46860 5528 47952 5556
rect 47946 5516 47952 5528
rect 48004 5516 48010 5568
rect 48608 5556 48636 5596
rect 48774 5584 48780 5596
rect 48832 5584 48838 5636
rect 50154 5556 50160 5568
rect 48608 5528 50160 5556
rect 50154 5516 50160 5528
rect 50212 5516 50218 5568
rect 50249 5559 50307 5565
rect 50249 5525 50261 5559
rect 50295 5556 50307 5559
rect 51074 5556 51080 5568
rect 50295 5528 51080 5556
rect 50295 5525 50307 5528
rect 50249 5519 50307 5525
rect 51074 5516 51080 5528
rect 51132 5516 51138 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 7098 5352 7104 5364
rect 1728 5324 7104 5352
rect 1728 5312 1734 5324
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 8352 5324 10701 5352
rect 8352 5312 8358 5324
rect 10689 5321 10701 5324
rect 10735 5321 10747 5355
rect 10689 5315 10747 5321
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14458 5352 14464 5364
rect 14323 5324 14464 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 17770 5312 17776 5364
rect 17828 5352 17834 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 17828 5324 18061 5352
rect 17828 5312 17834 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 21266 5352 21272 5364
rect 20864 5324 21272 5352
rect 20864 5312 20870 5324
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 24854 5352 24860 5364
rect 24815 5324 24860 5352
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 34422 5352 34428 5364
rect 33244 5324 34428 5352
rect 1854 5284 1860 5296
rect 1815 5256 1860 5284
rect 1854 5244 1860 5256
rect 1912 5244 1918 5296
rect 10042 5284 10048 5296
rect 2700 5256 10048 5284
rect 2700 5225 2728 5256
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 13164 5287 13222 5293
rect 10376 5256 10824 5284
rect 10376 5244 10382 5256
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 2685 5179 2743 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5040 5188 5549 5216
rect 5040 5176 5046 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7098 5216 7104 5228
rect 6972 5188 7017 5216
rect 7059 5188 7104 5216
rect 6972 5176 6978 5188
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10796 5225 10824 5256
rect 13164 5253 13176 5287
rect 13210 5284 13222 5287
rect 14090 5284 14096 5296
rect 13210 5256 14096 5284
rect 13210 5253 13222 5256
rect 13164 5247 13222 5253
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 20156 5287 20214 5293
rect 20156 5253 20168 5287
rect 20202 5284 20214 5287
rect 21818 5284 21824 5296
rect 20202 5256 21824 5284
rect 20202 5253 20214 5256
rect 20156 5247 20214 5253
rect 21818 5244 21824 5256
rect 21876 5244 21882 5296
rect 33042 5284 33048 5296
rect 25976 5256 33048 5284
rect 25976 5228 26004 5256
rect 33042 5244 33048 5256
rect 33100 5244 33106 5296
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 15378 5216 15384 5228
rect 10781 5179 10839 5185
rect 11164 5188 15384 5216
rect 2133 5151 2191 5157
rect 2133 5117 2145 5151
rect 2179 5148 2191 5151
rect 11164 5148 11192 5188
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 16925 5219 16983 5225
rect 16925 5216 16937 5219
rect 16816 5188 16937 5216
rect 16816 5176 16822 5188
rect 16925 5185 16937 5188
rect 16971 5185 16983 5219
rect 16925 5179 16983 5185
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19392 5188 19901 5216
rect 19392 5176 19398 5188
rect 19889 5185 19901 5188
rect 19935 5216 19947 5219
rect 20530 5216 20536 5228
rect 19935 5188 20536 5216
rect 19935 5185 19947 5188
rect 19889 5179 19947 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 24210 5216 24216 5228
rect 24171 5188 24216 5216
rect 24210 5176 24216 5188
rect 24268 5176 24274 5228
rect 24397 5219 24455 5225
rect 24397 5185 24409 5219
rect 24443 5216 24455 5219
rect 25041 5219 25099 5225
rect 25041 5216 25053 5219
rect 24443 5188 25053 5216
rect 24443 5185 24455 5188
rect 24397 5179 24455 5185
rect 25041 5185 25053 5188
rect 25087 5185 25099 5219
rect 25590 5216 25596 5228
rect 25551 5188 25596 5216
rect 25041 5179 25099 5185
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 25774 5216 25780 5228
rect 25735 5188 25780 5216
rect 25774 5176 25780 5188
rect 25832 5176 25838 5228
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26016 5188 26109 5216
rect 26016 5176 26022 5188
rect 26142 5176 26148 5228
rect 26200 5216 26206 5228
rect 27614 5216 27620 5228
rect 26200 5188 27620 5216
rect 26200 5176 26206 5188
rect 27614 5176 27620 5188
rect 27672 5176 27678 5228
rect 31297 5219 31355 5225
rect 31297 5185 31309 5219
rect 31343 5216 31355 5219
rect 33244 5216 33272 5324
rect 34422 5312 34428 5324
rect 34480 5312 34486 5364
rect 35986 5352 35992 5364
rect 35544 5324 35992 5352
rect 35342 5284 35348 5296
rect 34164 5256 35348 5284
rect 34164 5225 34192 5256
rect 35342 5244 35348 5256
rect 35400 5244 35406 5296
rect 35544 5293 35572 5324
rect 35986 5312 35992 5324
rect 36044 5312 36050 5364
rect 36078 5312 36084 5364
rect 36136 5352 36142 5364
rect 40310 5352 40316 5364
rect 36136 5324 40316 5352
rect 36136 5312 36142 5324
rect 40310 5312 40316 5324
rect 40368 5312 40374 5364
rect 35520 5287 35578 5293
rect 35520 5253 35532 5287
rect 35566 5253 35578 5287
rect 35520 5247 35578 5253
rect 39108 5287 39166 5293
rect 39108 5253 39120 5287
rect 39154 5284 39166 5287
rect 39206 5284 39212 5296
rect 39154 5256 39212 5284
rect 39154 5253 39166 5256
rect 39108 5247 39166 5253
rect 39206 5244 39212 5256
rect 39264 5244 39270 5296
rect 40218 5244 40224 5296
rect 40276 5284 40282 5296
rect 41046 5284 41052 5296
rect 40276 5256 41052 5284
rect 40276 5244 40282 5256
rect 41046 5244 41052 5256
rect 41104 5244 41110 5296
rect 51074 5293 51080 5296
rect 51068 5284 51080 5293
rect 51035 5256 51080 5284
rect 51068 5247 51080 5256
rect 51074 5244 51080 5247
rect 51132 5244 51138 5296
rect 31343 5188 33272 5216
rect 34057 5219 34115 5225
rect 31343 5185 31355 5188
rect 31297 5179 31355 5185
rect 34057 5185 34069 5219
rect 34103 5185 34115 5219
rect 34057 5179 34115 5185
rect 34149 5219 34207 5225
rect 34149 5185 34161 5219
rect 34195 5185 34207 5219
rect 34149 5179 34207 5185
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 2179 5120 11192 5148
rect 12406 5120 12909 5148
rect 2179 5117 2191 5120
rect 2133 5111 2191 5117
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 4065 5083 4123 5089
rect 4065 5080 4077 5083
rect 2832 5052 4077 5080
rect 2832 5040 2838 5052
rect 4065 5049 4077 5052
rect 4111 5049 4123 5083
rect 4065 5043 4123 5049
rect 9582 5040 9588 5092
rect 9640 5080 9646 5092
rect 10134 5080 10140 5092
rect 9640 5052 10140 5080
rect 9640 5040 9646 5052
rect 10134 5040 10140 5052
rect 10192 5080 10198 5092
rect 12406 5080 12434 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 10192 5052 12434 5080
rect 10192 5040 10198 5052
rect 2866 5012 2872 5024
rect 2827 4984 2872 5012
rect 2866 4972 2872 4984
rect 2924 4972 2930 5024
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 3878 5012 3884 5024
rect 3467 4984 3884 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 4709 5015 4767 5021
rect 4709 4981 4721 5015
rect 4755 5012 4767 5015
rect 5258 5012 5264 5024
rect 4755 4984 5264 5012
rect 4755 4981 4767 4984
rect 4709 4975 4767 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5353 5015 5411 5021
rect 5353 4981 5365 5015
rect 5399 5012 5411 5015
rect 6730 5012 6736 5024
rect 5399 4984 6736 5012
rect 5399 4981 5411 4984
rect 5353 4975 5411 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10410 5012 10416 5024
rect 10367 4984 10416 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 12912 5012 12940 5111
rect 15470 5012 15476 5024
rect 12912 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 5012 15534 5024
rect 16684 5012 16712 5111
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 24029 5151 24087 5157
rect 24029 5148 24041 5151
rect 22520 5120 24041 5148
rect 22520 5108 22526 5120
rect 24029 5117 24041 5120
rect 24075 5148 24087 5151
rect 24486 5148 24492 5160
rect 24075 5120 24492 5148
rect 24075 5117 24087 5120
rect 24029 5111 24087 5117
rect 24486 5108 24492 5120
rect 24544 5108 24550 5160
rect 25866 5148 25872 5160
rect 25827 5120 25872 5148
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 24762 5040 24768 5092
rect 24820 5080 24826 5092
rect 31312 5080 31340 5179
rect 33042 5108 33048 5160
rect 33100 5148 33106 5160
rect 34072 5148 34100 5179
rect 34330 5176 34336 5228
rect 34388 5216 34394 5228
rect 34425 5219 34483 5225
rect 34425 5216 34437 5219
rect 34388 5188 34437 5216
rect 34388 5176 34394 5188
rect 34425 5185 34437 5188
rect 34471 5185 34483 5219
rect 34425 5179 34483 5185
rect 35253 5219 35311 5225
rect 35253 5185 35265 5219
rect 35299 5216 35311 5219
rect 35299 5188 37964 5216
rect 35299 5185 35311 5188
rect 35253 5179 35311 5185
rect 37936 5160 37964 5188
rect 48590 5176 48596 5228
rect 48648 5216 48654 5228
rect 50801 5219 50859 5225
rect 50801 5216 50813 5219
rect 48648 5188 50813 5216
rect 48648 5176 48654 5188
rect 50801 5185 50813 5188
rect 50847 5185 50859 5219
rect 50801 5179 50859 5185
rect 33100 5120 34100 5148
rect 33100 5108 33106 5120
rect 37918 5108 37924 5160
rect 37976 5148 37982 5160
rect 38841 5151 38899 5157
rect 38841 5148 38853 5151
rect 37976 5120 38853 5148
rect 37976 5108 37982 5120
rect 38841 5117 38853 5120
rect 38887 5117 38899 5151
rect 38841 5111 38899 5117
rect 24820 5052 31340 5080
rect 31481 5083 31539 5089
rect 24820 5040 24826 5052
rect 31481 5049 31493 5083
rect 31527 5080 31539 5083
rect 35250 5080 35256 5092
rect 31527 5052 35256 5080
rect 31527 5049 31539 5052
rect 31481 5043 31539 5049
rect 15528 4984 16712 5012
rect 15528 4972 15534 4984
rect 30466 4972 30472 5024
rect 30524 5012 30530 5024
rect 31496 5012 31524 5043
rect 35250 5040 35256 5052
rect 35308 5040 35314 5092
rect 30524 4984 31524 5012
rect 30524 4972 30530 4984
rect 33502 4972 33508 5024
rect 33560 5012 33566 5024
rect 33873 5015 33931 5021
rect 33873 5012 33885 5015
rect 33560 4984 33885 5012
rect 33560 4972 33566 4984
rect 33873 4981 33885 4984
rect 33919 4981 33931 5015
rect 33873 4975 33931 4981
rect 34238 4972 34244 5024
rect 34296 5012 34302 5024
rect 34333 5015 34391 5021
rect 34333 5012 34345 5015
rect 34296 4984 34345 5012
rect 34296 4972 34302 4984
rect 34333 4981 34345 4984
rect 34379 4981 34391 5015
rect 34333 4975 34391 4981
rect 35894 4972 35900 5024
rect 35952 5012 35958 5024
rect 36633 5015 36691 5021
rect 36633 5012 36645 5015
rect 35952 4984 36645 5012
rect 35952 4972 35958 4984
rect 36633 4981 36645 4984
rect 36679 4981 36691 5015
rect 38856 5012 38884 5111
rect 41966 5080 41972 5092
rect 39776 5052 41972 5080
rect 39776 5012 39804 5052
rect 41966 5040 41972 5052
rect 42024 5040 42030 5092
rect 38856 4984 39804 5012
rect 36633 4975 36691 4981
rect 40126 4972 40132 5024
rect 40184 5012 40190 5024
rect 40221 5015 40279 5021
rect 40221 5012 40233 5015
rect 40184 4984 40233 5012
rect 40184 4972 40190 4984
rect 40221 4981 40233 4984
rect 40267 4981 40279 5015
rect 40221 4975 40279 4981
rect 48958 4972 48964 5024
rect 49016 5012 49022 5024
rect 52178 5012 52184 5024
rect 49016 4984 52184 5012
rect 49016 4972 49022 4984
rect 52178 4972 52184 4984
rect 52236 4972 52242 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 7466 4808 7472 4820
rect 2424 4780 7328 4808
rect 7427 4780 7472 4808
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2424 4613 2452 4780
rect 5166 4740 5172 4752
rect 5127 4712 5172 4740
rect 5166 4700 5172 4712
rect 5224 4700 5230 4752
rect 7300 4740 7328 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 11517 4811 11575 4817
rect 11517 4808 11529 4811
rect 10100 4780 11529 4808
rect 10100 4768 10106 4780
rect 11517 4777 11529 4780
rect 11563 4777 11575 4811
rect 11517 4771 11575 4777
rect 16669 4811 16727 4817
rect 16669 4777 16681 4811
rect 16715 4808 16727 4811
rect 16758 4808 16764 4820
rect 16715 4780 16764 4808
rect 16715 4777 16727 4780
rect 16669 4771 16727 4777
rect 16758 4768 16764 4780
rect 16816 4768 16822 4820
rect 24210 4768 24216 4820
rect 24268 4808 24274 4820
rect 25041 4811 25099 4817
rect 25041 4808 25053 4811
rect 24268 4780 25053 4808
rect 24268 4768 24274 4780
rect 25041 4777 25053 4780
rect 25087 4777 25099 4811
rect 30650 4808 30656 4820
rect 30611 4780 30656 4808
rect 25041 4771 25099 4777
rect 30650 4768 30656 4780
rect 30708 4768 30714 4820
rect 35526 4768 35532 4820
rect 35584 4768 35590 4820
rect 35986 4808 35992 4820
rect 35947 4780 35992 4808
rect 35986 4768 35992 4780
rect 36044 4768 36050 4820
rect 38654 4768 38660 4820
rect 38712 4808 38718 4820
rect 40405 4811 40463 4817
rect 40405 4808 40417 4811
rect 38712 4780 40417 4808
rect 38712 4768 38718 4780
rect 40405 4777 40417 4780
rect 40451 4777 40463 4811
rect 40405 4771 40463 4777
rect 48774 4768 48780 4820
rect 48832 4808 48838 4820
rect 49237 4811 49295 4817
rect 49237 4808 49249 4811
rect 48832 4780 49249 4808
rect 48832 4768 48838 4780
rect 49237 4777 49249 4780
rect 49283 4777 49295 4811
rect 49237 4771 49295 4777
rect 9582 4740 9588 4752
rect 7300 4712 9588 4740
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 19518 4740 19524 4752
rect 15948 4712 19524 4740
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4573 2467 4607
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 2409 4567 2467 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 4045 4607 4103 4613
rect 4045 4604 4057 4607
rect 3936 4576 4057 4604
rect 3936 4564 3942 4576
rect 4045 4573 4057 4576
rect 4091 4573 4103 4607
rect 4045 4567 4103 4573
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 6086 4604 6092 4616
rect 5592 4576 6092 4604
rect 5592 4564 5598 4576
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6914 4604 6920 4616
rect 6196 4576 6920 4604
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 6196 4536 6224 4576
rect 6914 4564 6920 4576
rect 6972 4604 6978 4616
rect 7742 4604 7748 4616
rect 6972 4576 7748 4604
rect 6972 4564 6978 4576
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 7926 4604 7932 4616
rect 7887 4576 7932 4604
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 9766 4604 9772 4616
rect 8159 4576 9772 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10410 4613 10416 4616
rect 10404 4604 10416 4613
rect 10371 4576 10416 4604
rect 10404 4567 10416 4576
rect 10410 4564 10416 4567
rect 10468 4564 10474 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 15948 4613 15976 4712
rect 19518 4700 19524 4712
rect 19576 4700 19582 4752
rect 26050 4740 26056 4752
rect 24504 4712 26056 4740
rect 16390 4672 16396 4684
rect 16224 4644 16396 4672
rect 16224 4613 16252 4644
rect 16390 4632 16396 4644
rect 16448 4672 16454 4684
rect 22278 4672 22284 4684
rect 16448 4644 17172 4672
rect 16448 4632 16454 4644
rect 17144 4613 17172 4644
rect 17880 4644 22284 4672
rect 15933 4607 15991 4613
rect 15933 4604 15945 4607
rect 13688 4576 15945 4604
rect 13688 4564 13694 4576
rect 15933 4573 15945 4576
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4573 16267 4607
rect 16209 4567 16267 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 3752 4508 6224 4536
rect 6356 4539 6414 4545
rect 3752 4496 3758 4508
rect 6356 4505 6368 4539
rect 6402 4536 6414 4539
rect 6638 4536 6644 4548
rect 6402 4508 6644 4536
rect 6402 4505 6414 4508
rect 6356 4499 6414 4505
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 13538 4496 13544 4548
rect 13596 4536 13602 4548
rect 16117 4539 16175 4545
rect 13596 4508 16068 4536
rect 13596 4496 13602 4508
rect 1578 4428 1584 4480
rect 1636 4468 1642 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1636 4440 1869 4468
rect 1636 4428 1642 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 1857 4431 1915 4437
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 2958 4468 2964 4480
rect 2639 4440 2964 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 7098 4468 7104 4480
rect 5224 4440 7104 4468
rect 5224 4428 5230 4440
rect 7098 4428 7104 4440
rect 7156 4468 7162 4480
rect 7834 4468 7840 4480
rect 7156 4440 7840 4468
rect 7156 4428 7162 4440
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 15746 4468 15752 4480
rect 15707 4440 15752 4468
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16040 4468 16068 4508
rect 16117 4505 16129 4539
rect 16163 4536 16175 4539
rect 16574 4536 16580 4548
rect 16163 4508 16580 4536
rect 16163 4505 16175 4508
rect 16117 4499 16175 4505
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16868 4468 16896 4567
rect 17037 4539 17095 4545
rect 17037 4505 17049 4539
rect 17083 4536 17095 4539
rect 17770 4536 17776 4548
rect 17083 4508 17776 4536
rect 17083 4505 17095 4508
rect 17037 4499 17095 4505
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 17880 4468 17908 4644
rect 22278 4632 22284 4644
rect 22336 4672 22342 4684
rect 23290 4672 23296 4684
rect 22336 4644 23296 4672
rect 22336 4632 22342 4644
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 24504 4672 24532 4712
rect 26050 4700 26056 4712
rect 26108 4700 26114 4752
rect 28994 4700 29000 4752
rect 29052 4740 29058 4752
rect 31665 4743 31723 4749
rect 31665 4740 31677 4743
rect 29052 4712 31677 4740
rect 29052 4700 29058 4712
rect 31665 4709 31677 4712
rect 31711 4709 31723 4743
rect 31665 4703 31723 4709
rect 33226 4700 33232 4752
rect 33284 4740 33290 4752
rect 33870 4740 33876 4752
rect 33284 4712 33876 4740
rect 33284 4700 33290 4712
rect 33870 4700 33876 4712
rect 33928 4700 33934 4752
rect 34238 4672 34244 4684
rect 24412 4644 24532 4672
rect 24688 4644 34244 4672
rect 19337 4607 19395 4613
rect 19337 4573 19349 4607
rect 19383 4604 19395 4607
rect 20254 4604 20260 4616
rect 19383 4576 20260 4604
rect 19383 4573 19395 4576
rect 19337 4567 19395 4573
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 22646 4564 22652 4616
rect 22704 4604 22710 4616
rect 24412 4613 24440 4644
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 22704 4576 24409 4604
rect 22704 4564 22710 4576
rect 24397 4573 24409 4576
rect 24443 4573 24455 4607
rect 24397 4567 24455 4573
rect 24486 4564 24492 4616
rect 24544 4604 24550 4616
rect 24688 4613 24716 4644
rect 24673 4607 24731 4613
rect 24544 4576 24589 4604
rect 24544 4564 24550 4576
rect 24673 4573 24685 4607
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 24854 4564 24860 4616
rect 24912 4613 24918 4616
rect 24912 4604 24920 4613
rect 24912 4576 24957 4604
rect 24912 4567 24920 4576
rect 24912 4564 24918 4567
rect 25130 4564 25136 4616
rect 25188 4604 25194 4616
rect 26142 4604 26148 4616
rect 25188 4576 26148 4604
rect 25188 4564 25194 4576
rect 26142 4564 26148 4576
rect 26200 4564 26206 4616
rect 27816 4613 27844 4644
rect 34238 4632 34244 4644
rect 34296 4632 34302 4684
rect 35544 4681 35572 4768
rect 37458 4700 37464 4752
rect 37516 4740 37522 4752
rect 37829 4743 37887 4749
rect 37829 4740 37841 4743
rect 37516 4712 37841 4740
rect 37516 4700 37522 4712
rect 37829 4709 37841 4712
rect 37875 4740 37887 4743
rect 40310 4740 40316 4752
rect 37875 4712 40316 4740
rect 37875 4709 37887 4712
rect 37829 4703 37887 4709
rect 40310 4700 40316 4712
rect 40368 4740 40374 4752
rect 48866 4740 48872 4752
rect 40368 4712 48872 4740
rect 40368 4700 40374 4712
rect 48866 4700 48872 4712
rect 48924 4700 48930 4752
rect 35529 4675 35587 4681
rect 35529 4641 35541 4675
rect 35575 4641 35587 4675
rect 35529 4635 35587 4641
rect 36078 4632 36084 4684
rect 36136 4672 36142 4684
rect 39758 4672 39764 4684
rect 36136 4644 39764 4672
rect 36136 4632 36142 4644
rect 39758 4632 39764 4644
rect 39816 4632 39822 4684
rect 40034 4632 40040 4684
rect 40092 4672 40098 4684
rect 40092 4644 40264 4672
rect 40092 4632 40098 4644
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 29546 4564 29552 4616
rect 29604 4604 29610 4616
rect 30101 4607 30159 4613
rect 30101 4604 30113 4607
rect 29604 4576 30113 4604
rect 29604 4564 29610 4576
rect 30101 4573 30113 4576
rect 30147 4573 30159 4607
rect 30466 4604 30472 4616
rect 30427 4576 30472 4604
rect 30101 4567 30159 4573
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 31110 4604 31116 4616
rect 31071 4576 31116 4604
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 31481 4607 31539 4613
rect 31481 4573 31493 4607
rect 31527 4604 31539 4607
rect 31570 4604 31576 4616
rect 31527 4576 31576 4604
rect 31527 4573 31539 4576
rect 31481 4567 31539 4573
rect 31570 4564 31576 4576
rect 31628 4564 31634 4616
rect 33318 4604 33324 4616
rect 33279 4576 33324 4604
rect 33318 4564 33324 4576
rect 33376 4564 33382 4616
rect 33502 4604 33508 4616
rect 33463 4576 33508 4604
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 33686 4564 33692 4616
rect 33744 4604 33750 4616
rect 33744 4576 33789 4604
rect 33744 4564 33750 4576
rect 35250 4564 35256 4616
rect 35308 4564 35314 4616
rect 35434 4613 35440 4616
rect 35409 4607 35440 4613
rect 35409 4573 35421 4607
rect 35409 4567 35440 4573
rect 35434 4564 35440 4567
rect 35492 4564 35498 4616
rect 35710 4613 35716 4616
rect 35667 4607 35716 4613
rect 35667 4573 35679 4607
rect 35713 4573 35716 4607
rect 35667 4567 35716 4573
rect 35710 4564 35716 4567
rect 35768 4564 35774 4616
rect 35805 4607 35863 4613
rect 35805 4573 35817 4607
rect 35851 4604 35863 4607
rect 35894 4604 35900 4616
rect 35851 4576 35900 4604
rect 35851 4573 35863 4576
rect 35805 4567 35863 4573
rect 35894 4564 35900 4576
rect 35952 4564 35958 4616
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 37645 4607 37703 4613
rect 37645 4604 37657 4607
rect 37608 4576 37657 4604
rect 37608 4564 37614 4576
rect 37645 4573 37657 4576
rect 37691 4573 37703 4607
rect 39850 4604 39856 4616
rect 39811 4576 39856 4604
rect 37645 4567 37703 4573
rect 39850 4564 39856 4576
rect 39908 4564 39914 4616
rect 40126 4604 40132 4616
rect 40087 4576 40132 4604
rect 40126 4564 40132 4576
rect 40184 4564 40190 4616
rect 40236 4613 40264 4644
rect 40770 4632 40776 4684
rect 40828 4672 40834 4684
rect 45462 4672 45468 4684
rect 40828 4644 45468 4672
rect 40828 4632 40834 4644
rect 45462 4632 45468 4644
rect 45520 4672 45526 4684
rect 45649 4675 45707 4681
rect 45649 4672 45661 4675
rect 45520 4644 45661 4672
rect 45520 4632 45526 4644
rect 45649 4641 45661 4644
rect 45695 4641 45707 4675
rect 45649 4635 45707 4641
rect 46290 4632 46296 4684
rect 46348 4672 46354 4684
rect 47118 4672 47124 4684
rect 46348 4644 47124 4672
rect 46348 4632 46354 4644
rect 47118 4632 47124 4644
rect 47176 4672 47182 4684
rect 47486 4672 47492 4684
rect 47176 4644 47492 4672
rect 47176 4632 47182 4644
rect 47486 4632 47492 4644
rect 47544 4672 47550 4684
rect 48038 4672 48044 4684
rect 47544 4644 48044 4672
rect 47544 4632 47550 4644
rect 48038 4632 48044 4644
rect 48096 4632 48102 4684
rect 48516 4644 49096 4672
rect 40221 4607 40279 4613
rect 40221 4573 40233 4607
rect 40267 4604 40279 4607
rect 46845 4607 46903 4613
rect 46845 4604 46857 4607
rect 40267 4576 46857 4604
rect 40267 4573 40279 4576
rect 40221 4567 40279 4573
rect 46845 4573 46857 4576
rect 46891 4604 46903 4607
rect 48516 4604 48544 4644
rect 48682 4604 48688 4616
rect 46891 4576 48544 4604
rect 48643 4576 48688 4604
rect 46891 4573 46903 4576
rect 46845 4567 46903 4573
rect 48682 4564 48688 4576
rect 48740 4564 48746 4616
rect 48866 4604 48872 4616
rect 48827 4576 48872 4604
rect 48866 4564 48872 4576
rect 48924 4564 48930 4616
rect 49068 4613 49096 4644
rect 49053 4607 49111 4613
rect 49053 4573 49065 4607
rect 49099 4604 49111 4607
rect 49142 4604 49148 4616
rect 49099 4576 49148 4604
rect 49099 4573 49111 4576
rect 49053 4567 49111 4573
rect 49142 4564 49148 4576
rect 49200 4564 49206 4616
rect 19518 4536 19524 4548
rect 19479 4508 19524 4536
rect 19518 4496 19524 4508
rect 19576 4536 19582 4548
rect 20438 4536 20444 4548
rect 19576 4508 20444 4536
rect 19576 4496 19582 4508
rect 20438 4496 20444 4508
rect 20496 4496 20502 4548
rect 24302 4496 24308 4548
rect 24360 4536 24366 4548
rect 24765 4539 24823 4545
rect 24765 4536 24777 4539
rect 24360 4508 24777 4536
rect 24360 4496 24366 4508
rect 24765 4505 24777 4508
rect 24811 4536 24823 4539
rect 25866 4536 25872 4548
rect 24811 4508 25872 4536
rect 24811 4505 24823 4508
rect 24765 4499 24823 4505
rect 25866 4496 25872 4508
rect 25924 4496 25930 4548
rect 27982 4536 27988 4548
rect 27895 4508 27988 4536
rect 27982 4496 27988 4508
rect 28040 4536 28046 4548
rect 30190 4536 30196 4548
rect 28040 4508 30196 4536
rect 28040 4496 28046 4508
rect 30190 4496 30196 4508
rect 30248 4536 30254 4548
rect 30285 4539 30343 4545
rect 30285 4536 30297 4539
rect 30248 4508 30297 4536
rect 30248 4496 30254 4508
rect 30285 4505 30297 4508
rect 30331 4505 30343 4539
rect 30285 4499 30343 4505
rect 30377 4539 30435 4545
rect 30377 4505 30389 4539
rect 30423 4536 30435 4539
rect 30926 4536 30932 4548
rect 30423 4508 30932 4536
rect 30423 4505 30435 4508
rect 30377 4499 30435 4505
rect 30926 4496 30932 4508
rect 30984 4496 30990 4548
rect 31294 4536 31300 4548
rect 31255 4508 31300 4536
rect 31294 4496 31300 4508
rect 31352 4496 31358 4548
rect 31389 4539 31447 4545
rect 31389 4505 31401 4539
rect 31435 4536 31447 4539
rect 33134 4536 33140 4548
rect 31435 4508 33140 4536
rect 31435 4505 31447 4508
rect 31389 4499 31447 4505
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 33594 4536 33600 4548
rect 33555 4508 33600 4536
rect 33594 4496 33600 4508
rect 33652 4496 33658 4548
rect 16040 4440 17908 4468
rect 19426 4428 19432 4480
rect 19484 4468 19490 4480
rect 19705 4471 19763 4477
rect 19705 4468 19717 4471
rect 19484 4440 19717 4468
rect 19484 4428 19490 4440
rect 19705 4437 19717 4440
rect 19751 4437 19763 4471
rect 19705 4431 19763 4437
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 27706 4468 27712 4480
rect 22152 4440 27712 4468
rect 22152 4428 22158 4440
rect 27706 4428 27712 4440
rect 27764 4428 27770 4480
rect 31570 4428 31576 4480
rect 31628 4468 31634 4480
rect 33704 4468 33732 4564
rect 35253 4551 35265 4564
rect 35299 4551 35311 4564
rect 35253 4545 35311 4551
rect 40037 4539 40095 4545
rect 40037 4505 40049 4539
rect 40083 4536 40095 4539
rect 40310 4536 40316 4548
rect 40083 4508 40316 4536
rect 40083 4505 40095 4508
rect 40037 4499 40095 4505
rect 40310 4496 40316 4508
rect 40368 4496 40374 4548
rect 40957 4539 41015 4545
rect 40957 4505 40969 4539
rect 41003 4536 41015 4539
rect 45094 4536 45100 4548
rect 41003 4508 45100 4536
rect 41003 4505 41015 4508
rect 40957 4499 41015 4505
rect 45094 4496 45100 4508
rect 45152 4536 45158 4548
rect 45465 4539 45523 4545
rect 45465 4536 45477 4539
rect 45152 4508 45477 4536
rect 45152 4496 45158 4508
rect 45465 4505 45477 4508
rect 45511 4505 45523 4539
rect 45465 4499 45523 4505
rect 48314 4496 48320 4548
rect 48372 4536 48378 4548
rect 48958 4536 48964 4548
rect 48372 4508 48964 4536
rect 48372 4496 48378 4508
rect 48958 4496 48964 4508
rect 49016 4496 49022 4548
rect 31628 4440 33732 4468
rect 33873 4471 33931 4477
rect 31628 4428 31634 4440
rect 33873 4437 33885 4471
rect 33919 4468 33931 4471
rect 33962 4468 33968 4480
rect 33919 4440 33968 4468
rect 33919 4437 33931 4440
rect 33873 4431 33931 4437
rect 33962 4428 33968 4440
rect 34020 4428 34026 4480
rect 34238 4428 34244 4480
rect 34296 4468 34302 4480
rect 37550 4468 37556 4480
rect 34296 4440 37556 4468
rect 34296 4428 34302 4440
rect 37550 4428 37556 4440
rect 37608 4428 37614 4480
rect 37734 4428 37740 4480
rect 37792 4468 37798 4480
rect 41049 4471 41107 4477
rect 41049 4468 41061 4471
rect 37792 4440 41061 4468
rect 37792 4428 37798 4440
rect 41049 4437 41061 4440
rect 41095 4468 41107 4471
rect 41230 4468 41236 4480
rect 41095 4440 41236 4468
rect 41095 4437 41107 4440
rect 41049 4431 41107 4437
rect 41230 4428 41236 4440
rect 41288 4428 41294 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3326 4264 3332 4276
rect 3239 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3973 4267 4031 4273
rect 3973 4233 3985 4267
rect 4019 4233 4031 4267
rect 3973 4227 4031 4233
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4233 5227 4267
rect 6638 4264 6644 4276
rect 6599 4236 6644 4264
rect 5169 4227 5227 4233
rect 2216 4131 2274 4137
rect 2216 4097 2228 4131
rect 2262 4128 2274 4131
rect 2774 4128 2780 4140
rect 2262 4100 2780 4128
rect 2262 4097 2274 4100
rect 2216 4091 2274 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3344 4128 3372 4224
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 3988 4196 4016 4227
rect 3936 4168 4016 4196
rect 3936 4156 3942 4168
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 4982 4196 4988 4208
rect 4212 4168 4988 4196
rect 4212 4156 4218 4168
rect 4982 4156 4988 4168
rect 5040 4156 5046 4208
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5184 4196 5212 4227
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 7926 4264 7932 4276
rect 6788 4236 6833 4264
rect 7887 4236 7932 4264
rect 6788 4224 6794 4236
rect 7926 4224 7932 4236
rect 7984 4224 7990 4276
rect 14921 4267 14979 4273
rect 14921 4233 14933 4267
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 5442 4196 5448 4208
rect 5132 4168 5212 4196
rect 5276 4168 5448 4196
rect 5132 4156 5138 4168
rect 3694 4128 3700 4140
rect 3344 4100 3700 4128
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 5276 4128 5304 4168
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 6656 4168 6960 4196
rect 3835 4100 5304 4128
rect 5353 4131 5411 4137
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5534 4128 5540 4140
rect 5399 4100 5540 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6546 4128 6552 4140
rect 6411 4100 6552 4128
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 6546 4088 6552 4100
rect 6604 4128 6610 4140
rect 6656 4128 6684 4168
rect 6822 4128 6828 4140
rect 6604 4100 6684 4128
rect 6783 4100 6828 4128
rect 6604 4088 6610 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6932 4128 6960 4168
rect 7576 4168 7788 4196
rect 7576 4128 7604 4168
rect 6932 4100 7604 4128
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7760 4128 7788 4168
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 9364 4168 9720 4196
rect 9364 4156 9370 4168
rect 8386 4128 8392 4140
rect 7760 4100 8392 4128
rect 7653 4091 7711 4097
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 6638 4060 6644 4072
rect 3016 4032 6644 4060
rect 3016 4020 3022 4032
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 7668 4060 7696 4091
rect 7944 4069 7972 4100
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9582 4128 9588 4140
rect 9543 4100 9588 4128
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 9692 4128 9720 4168
rect 10336 4168 10824 4196
rect 10336 4128 10364 4168
rect 9692 4100 10364 4128
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10468 4100 10701 4128
rect 10468 4088 10474 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10796 4128 10824 4168
rect 12526 4156 12532 4208
rect 12584 4156 12590 4208
rect 13814 4156 13820 4208
rect 13872 4196 13878 4208
rect 13909 4199 13967 4205
rect 13909 4196 13921 4199
rect 13872 4168 13921 4196
rect 13872 4156 13878 4168
rect 13909 4165 13921 4168
rect 13955 4165 13967 4199
rect 13909 4159 13967 4165
rect 12544 4128 12572 4156
rect 10796 4100 12572 4128
rect 12713 4131 12771 4137
rect 10689 4091 10747 4097
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 12986 4128 12992 4140
rect 12759 4100 12992 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 6788 4032 7696 4060
rect 7929 4063 7987 4069
rect 6788 4020 6794 4032
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 12529 4063 12587 4069
rect 12529 4060 12541 4063
rect 8076 4032 12541 4060
rect 8076 4020 8082 4032
rect 12529 4029 12541 4032
rect 12575 4029 12587 4063
rect 14936 4060 14964 4227
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 24486 4264 24492 4276
rect 20220 4236 24492 4264
rect 20220 4224 20226 4236
rect 24486 4224 24492 4236
rect 24544 4224 24550 4276
rect 25774 4264 25780 4276
rect 25608 4236 25780 4264
rect 15010 4156 15016 4208
rect 15068 4196 15074 4208
rect 15068 4168 15240 4196
rect 15068 4156 15074 4168
rect 15102 4128 15108 4140
rect 15063 4100 15108 4128
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15212 4128 15240 4168
rect 16132 4168 16988 4196
rect 16132 4128 16160 4168
rect 15212 4100 16160 4128
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16264 4100 16865 4128
rect 16264 4088 16270 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16960 4128 16988 4168
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 25608 4196 25636 4236
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 31294 4224 31300 4276
rect 31352 4264 31358 4276
rect 31389 4267 31447 4273
rect 31389 4264 31401 4267
rect 31352 4236 31401 4264
rect 31352 4224 31358 4236
rect 31389 4233 31401 4236
rect 31435 4233 31447 4267
rect 31389 4227 31447 4233
rect 33042 4224 33048 4276
rect 33100 4264 33106 4276
rect 37458 4264 37464 4276
rect 33100 4236 37464 4264
rect 33100 4224 33106 4236
rect 37458 4224 37464 4236
rect 37516 4224 37522 4276
rect 41046 4224 41052 4276
rect 41104 4264 41110 4276
rect 43806 4264 43812 4276
rect 41104 4236 41736 4264
rect 43767 4236 43812 4264
rect 41104 4224 41110 4236
rect 29086 4196 29092 4208
rect 24912 4168 25636 4196
rect 24912 4156 24918 4168
rect 19058 4128 19064 4140
rect 16960 4100 19064 4128
rect 16853 4091 16911 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19426 4128 19432 4140
rect 19199 4100 19432 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 23290 4128 23296 4140
rect 22695 4100 23296 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 23624 4100 23857 4128
rect 23624 4088 23630 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 24394 4088 24400 4140
rect 24452 4128 24458 4140
rect 25409 4131 25467 4137
rect 25409 4128 25421 4131
rect 24452 4100 25421 4128
rect 24452 4088 24458 4100
rect 25409 4097 25421 4100
rect 25455 4128 25467 4131
rect 25498 4128 25504 4140
rect 25455 4100 25504 4128
rect 25455 4097 25467 4100
rect 25409 4091 25467 4097
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 25608 4137 25636 4168
rect 28276 4168 29092 4196
rect 25593 4131 25651 4137
rect 25593 4097 25605 4131
rect 25639 4097 25651 4131
rect 25593 4091 25651 4097
rect 25777 4131 25835 4137
rect 25777 4097 25789 4131
rect 25823 4128 25835 4131
rect 25866 4128 25872 4140
rect 25823 4100 25872 4128
rect 25823 4097 25835 4100
rect 25777 4091 25835 4097
rect 25866 4088 25872 4100
rect 25924 4088 25930 4140
rect 28276 4137 28304 4168
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 30944 4168 31156 4196
rect 25961 4131 26019 4137
rect 25961 4097 25973 4131
rect 26007 4097 26019 4131
rect 25961 4091 26019 4097
rect 28261 4131 28319 4137
rect 28261 4097 28273 4131
rect 28307 4097 28319 4131
rect 28261 4091 28319 4097
rect 28528 4131 28586 4137
rect 28528 4097 28540 4131
rect 28574 4128 28586 4131
rect 28994 4128 29000 4140
rect 28574 4100 29000 4128
rect 28574 4097 28586 4100
rect 28528 4091 28586 4097
rect 22370 4060 22376 4072
rect 14936 4032 22376 4060
rect 12529 4023 12587 4029
rect 22370 4020 22376 4032
rect 22428 4020 22434 4072
rect 22462 4020 22468 4072
rect 22520 4060 22526 4072
rect 22520 4032 22565 4060
rect 22520 4020 22526 4032
rect 23014 4020 23020 4072
rect 23072 4060 23078 4072
rect 25685 4063 25743 4069
rect 25685 4060 25697 4063
rect 23072 4032 25697 4060
rect 23072 4020 23078 4032
rect 25685 4029 25697 4032
rect 25731 4029 25743 4063
rect 25685 4023 25743 4029
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 3292 3964 5028 3992
rect 3292 3952 3298 3964
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 2188 3896 4721 3924
rect 2188 3884 2194 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 5000 3924 5028 3964
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 5132 3964 8401 3992
rect 5132 3952 5138 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 10134 3992 10140 4004
rect 8389 3955 8447 3961
rect 8496 3964 10140 3992
rect 6730 3924 6736 3936
rect 5000 3896 6736 3924
rect 4709 3887 4767 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 8018 3924 8024 3936
rect 7791 3896 8024 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8496 3924 8524 3964
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 10505 3995 10563 4001
rect 10505 3961 10517 3995
rect 10551 3992 10563 3995
rect 10594 3992 10600 4004
rect 10551 3964 10600 3992
rect 10551 3961 10563 3964
rect 10505 3955 10563 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 22094 3992 22100 4004
rect 10836 3964 22100 3992
rect 10836 3952 10842 3964
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 22186 3952 22192 4004
rect 22244 3992 22250 4004
rect 23658 3992 23664 4004
rect 22244 3964 23520 3992
rect 23619 3964 23664 3992
rect 22244 3952 22250 3964
rect 9674 3924 9680 3936
rect 8168 3896 8524 3924
rect 9635 3896 9680 3924
rect 8168 3884 8174 3896
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 11330 3924 11336 3936
rect 9824 3896 11336 3924
rect 9824 3884 9830 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 16022 3924 16028 3936
rect 12943 3896 16028 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 18966 3924 18972 3936
rect 18927 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 20254 3924 20260 3936
rect 19116 3896 20260 3924
rect 19116 3884 19122 3896
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 22833 3927 22891 3933
rect 22833 3924 22845 3927
rect 20404 3896 22845 3924
rect 20404 3884 20410 3896
rect 22833 3893 22845 3896
rect 22879 3893 22891 3927
rect 23492 3924 23520 3964
rect 23658 3952 23664 3964
rect 23716 3952 23722 4004
rect 25976 3936 26004 4091
rect 28994 4088 29000 4100
rect 29052 4088 29058 4140
rect 30282 4088 30288 4140
rect 30340 4128 30346 4140
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30340 4100 30849 4128
rect 30340 4088 30346 4100
rect 30837 4097 30849 4100
rect 30883 4097 30895 4131
rect 30837 4091 30895 4097
rect 29546 4020 29552 4072
rect 29604 4060 29610 4072
rect 30944 4060 30972 4168
rect 31128 4137 31156 4168
rect 36078 4156 36084 4208
rect 36136 4196 36142 4208
rect 40770 4196 40776 4208
rect 36136 4168 40776 4196
rect 36136 4156 36142 4168
rect 31021 4131 31079 4137
rect 31021 4097 31033 4131
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 31113 4131 31171 4137
rect 31113 4097 31125 4131
rect 31159 4097 31171 4131
rect 31113 4091 31171 4097
rect 31205 4131 31263 4137
rect 31205 4097 31217 4131
rect 31251 4128 31263 4131
rect 31938 4128 31944 4140
rect 31251 4100 31944 4128
rect 31251 4097 31263 4100
rect 31205 4091 31263 4097
rect 29604 4032 30972 4060
rect 31036 4060 31064 4091
rect 31938 4088 31944 4100
rect 31996 4088 32002 4140
rect 32122 4088 32128 4140
rect 32180 4128 32186 4140
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 32180 4100 32321 4128
rect 32180 4088 32186 4100
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 33778 4088 33784 4140
rect 33836 4128 33842 4140
rect 37461 4131 37519 4137
rect 33836 4100 37412 4128
rect 33836 4088 33842 4100
rect 33042 4060 33048 4072
rect 31036 4032 33048 4060
rect 29604 4020 29610 4032
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 35894 4020 35900 4072
rect 35952 4060 35958 4072
rect 37277 4063 37335 4069
rect 37277 4060 37289 4063
rect 35952 4032 37289 4060
rect 35952 4020 35958 4032
rect 37277 4029 37289 4032
rect 37323 4029 37335 4063
rect 37384 4060 37412 4100
rect 37461 4097 37473 4131
rect 37507 4128 37519 4131
rect 37826 4128 37832 4140
rect 37507 4100 37832 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 38304 4137 38332 4168
rect 40770 4156 40776 4168
rect 40828 4156 40834 4208
rect 38289 4131 38347 4137
rect 38289 4097 38301 4131
rect 38335 4097 38347 4131
rect 38289 4091 38347 4097
rect 38378 4088 38384 4140
rect 38436 4137 38442 4140
rect 38436 4131 38485 4137
rect 38436 4097 38439 4131
rect 38473 4097 38485 4131
rect 38562 4128 38568 4140
rect 38523 4100 38568 4128
rect 38436 4091 38485 4097
rect 38436 4088 38442 4091
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 38746 4137 38752 4140
rect 38703 4131 38752 4137
rect 38703 4097 38715 4131
rect 38749 4097 38752 4131
rect 38703 4091 38752 4097
rect 38746 4088 38752 4091
rect 38804 4088 38810 4140
rect 40405 4131 40463 4137
rect 40405 4097 40417 4131
rect 40451 4128 40463 4131
rect 41046 4128 41052 4140
rect 40451 4100 41052 4128
rect 40451 4097 40463 4100
rect 40405 4091 40463 4097
rect 41046 4088 41052 4100
rect 41104 4088 41110 4140
rect 41141 4131 41199 4137
rect 41141 4097 41153 4131
rect 41187 4128 41199 4131
rect 41230 4128 41236 4140
rect 41187 4100 41236 4128
rect 41187 4097 41199 4100
rect 41141 4091 41199 4097
rect 41230 4088 41236 4100
rect 41288 4088 41294 4140
rect 41325 4131 41383 4137
rect 41325 4097 41337 4131
rect 41371 4097 41383 4131
rect 41325 4091 41383 4097
rect 41417 4131 41475 4137
rect 41417 4097 41429 4131
rect 41463 4097 41475 4131
rect 41417 4091 41475 4097
rect 41533 4131 41591 4137
rect 41533 4097 41545 4131
rect 41579 4128 41591 4131
rect 41708 4128 41736 4236
rect 43806 4224 43812 4236
rect 43864 4224 43870 4276
rect 45462 4224 45468 4276
rect 45520 4264 45526 4276
rect 45520 4236 46520 4264
rect 45520 4224 45526 4236
rect 45649 4199 45707 4205
rect 45649 4165 45661 4199
rect 45695 4196 45707 4199
rect 46382 4196 46388 4208
rect 45695 4168 46388 4196
rect 45695 4165 45707 4168
rect 45649 4159 45707 4165
rect 46382 4156 46388 4168
rect 46440 4156 46446 4208
rect 42685 4131 42743 4137
rect 42685 4128 42697 4131
rect 41579 4100 41736 4128
rect 41892 4100 42697 4128
rect 41579 4097 41591 4100
rect 41533 4091 41591 4097
rect 37384 4032 41184 4060
rect 37277 4023 37335 4029
rect 33778 3992 33784 4004
rect 29472 3964 33784 3992
rect 25958 3924 25964 3936
rect 23492 3896 25964 3924
rect 22833 3887 22891 3893
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 26145 3927 26203 3933
rect 26145 3893 26157 3927
rect 26191 3924 26203 3927
rect 26418 3924 26424 3936
rect 26191 3896 26424 3924
rect 26191 3893 26203 3896
rect 26145 3887 26203 3893
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 26878 3884 26884 3936
rect 26936 3924 26942 3936
rect 29472 3924 29500 3964
rect 33778 3952 33784 3964
rect 33836 3952 33842 4004
rect 35802 3952 35808 4004
rect 35860 3992 35866 4004
rect 36630 3992 36636 4004
rect 35860 3964 36636 3992
rect 35860 3952 35866 3964
rect 36630 3952 36636 3964
rect 36688 3952 36694 4004
rect 38746 3952 38752 4004
rect 38804 3992 38810 4004
rect 40862 3992 40868 4004
rect 38804 3964 40868 3992
rect 38804 3952 38810 3964
rect 40862 3952 40868 3964
rect 40920 3952 40926 4004
rect 26936 3896 29500 3924
rect 26936 3884 26942 3896
rect 29546 3884 29552 3936
rect 29604 3924 29610 3936
rect 29641 3927 29699 3933
rect 29641 3924 29653 3927
rect 29604 3896 29653 3924
rect 29604 3884 29610 3896
rect 29641 3893 29653 3896
rect 29687 3893 29699 3927
rect 29641 3887 29699 3893
rect 30190 3884 30196 3936
rect 30248 3924 30254 3936
rect 32122 3924 32128 3936
rect 30248 3896 32128 3924
rect 30248 3884 30254 3896
rect 32122 3884 32128 3896
rect 32180 3884 32186 3936
rect 32490 3924 32496 3936
rect 32451 3896 32496 3924
rect 32490 3884 32496 3896
rect 32548 3884 32554 3936
rect 32582 3884 32588 3936
rect 32640 3924 32646 3936
rect 35342 3924 35348 3936
rect 32640 3896 35348 3924
rect 32640 3884 32646 3896
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 36446 3884 36452 3936
rect 36504 3924 36510 3936
rect 37645 3927 37703 3933
rect 37645 3924 37657 3927
rect 36504 3896 37657 3924
rect 36504 3884 36510 3896
rect 37645 3893 37657 3896
rect 37691 3893 37703 3927
rect 38838 3924 38844 3936
rect 38799 3896 38844 3924
rect 37645 3887 37703 3893
rect 38838 3884 38844 3896
rect 38896 3884 38902 3936
rect 40589 3927 40647 3933
rect 40589 3893 40601 3927
rect 40635 3924 40647 3927
rect 40954 3924 40960 3936
rect 40635 3896 40960 3924
rect 40635 3893 40647 3896
rect 40589 3887 40647 3893
rect 40954 3884 40960 3896
rect 41012 3884 41018 3936
rect 41156 3924 41184 4032
rect 41340 4004 41368 4091
rect 41432 4004 41460 4091
rect 41322 3952 41328 4004
rect 41380 3952 41386 4004
rect 41414 3952 41420 4004
rect 41472 3952 41478 4004
rect 41693 3995 41751 4001
rect 41693 3961 41705 3995
rect 41739 3992 41751 3995
rect 41892 3992 41920 4100
rect 42685 4097 42697 4100
rect 42731 4097 42743 4131
rect 45462 4128 45468 4140
rect 45423 4100 45468 4128
rect 42685 4091 42743 4097
rect 45462 4088 45468 4100
rect 45520 4088 45526 4140
rect 45738 4128 45744 4140
rect 45699 4100 45744 4128
rect 45738 4088 45744 4100
rect 45796 4088 45802 4140
rect 45830 4088 45836 4140
rect 45888 4128 45894 4140
rect 46492 4137 46520 4236
rect 48866 4224 48872 4276
rect 48924 4224 48930 4276
rect 46753 4199 46811 4205
rect 46753 4196 46765 4199
rect 46584 4168 46765 4196
rect 46477 4131 46535 4137
rect 45888 4100 45933 4128
rect 45888 4088 45894 4100
rect 46477 4097 46489 4131
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 41966 4020 41972 4072
rect 42024 4060 42030 4072
rect 42426 4060 42432 4072
rect 42024 4032 42432 4060
rect 42024 4020 42030 4032
rect 42426 4020 42432 4032
rect 42484 4020 42490 4072
rect 46584 4060 46612 4168
rect 46753 4165 46765 4168
rect 46799 4165 46811 4199
rect 46753 4159 46811 4165
rect 47026 4156 47032 4208
rect 47084 4196 47090 4208
rect 47765 4199 47823 4205
rect 47765 4196 47777 4199
rect 47084 4168 47777 4196
rect 47084 4156 47090 4168
rect 47765 4165 47777 4168
rect 47811 4165 47823 4199
rect 48682 4196 48688 4208
rect 47765 4159 47823 4165
rect 47872 4168 48688 4196
rect 46661 4131 46719 4137
rect 46661 4097 46673 4131
rect 46707 4097 46719 4131
rect 46842 4128 46848 4140
rect 46803 4100 46848 4128
rect 46661 4091 46719 4097
rect 45872 4032 46612 4060
rect 46676 4060 46704 4091
rect 46842 4088 46848 4100
rect 46900 4088 46906 4140
rect 47578 4128 47584 4140
rect 47539 4100 47584 4128
rect 47578 4088 47584 4100
rect 47636 4088 47642 4140
rect 47872 4137 47900 4168
rect 48682 4156 48688 4168
rect 48740 4156 48746 4208
rect 48884 4196 48912 4224
rect 48961 4199 49019 4205
rect 48961 4196 48973 4199
rect 48884 4168 48973 4196
rect 48961 4165 48973 4168
rect 49007 4165 49019 4199
rect 48961 4159 49019 4165
rect 47857 4131 47915 4137
rect 47857 4097 47869 4131
rect 47903 4097 47915 4131
rect 47857 4091 47915 4097
rect 47949 4131 48007 4137
rect 47949 4097 47961 4131
rect 47995 4128 48007 4131
rect 48038 4128 48044 4140
rect 47995 4100 48044 4128
rect 47995 4097 48007 4100
rect 47949 4091 48007 4097
rect 48038 4088 48044 4100
rect 48096 4088 48102 4140
rect 48774 4088 48780 4140
rect 48832 4137 48838 4140
rect 48832 4131 48855 4137
rect 48843 4097 48855 4131
rect 49050 4128 49056 4140
rect 49011 4100 49056 4128
rect 48832 4091 48855 4097
rect 48832 4088 48838 4091
rect 49050 4088 49056 4100
rect 49108 4088 49114 4140
rect 49142 4088 49148 4140
rect 49200 4128 49206 4140
rect 49200 4100 49245 4128
rect 49200 4088 49206 4100
rect 46676 4032 48176 4060
rect 41739 3964 41920 3992
rect 41739 3961 41751 3964
rect 41693 3955 41751 3961
rect 45872 3924 45900 4032
rect 46017 3995 46075 4001
rect 46017 3961 46029 3995
rect 46063 3992 46075 3995
rect 48038 3992 48044 4004
rect 46063 3964 48044 3992
rect 46063 3961 46075 3964
rect 46017 3955 46075 3961
rect 48038 3952 48044 3964
rect 48096 3952 48102 4004
rect 48148 4001 48176 4032
rect 48133 3995 48191 4001
rect 48133 3961 48145 3995
rect 48179 3961 48191 3995
rect 49326 3992 49332 4004
rect 49287 3964 49332 3992
rect 48133 3955 48191 3961
rect 49326 3952 49332 3964
rect 49384 3952 49390 4004
rect 47026 3924 47032 3936
rect 41156 3896 45900 3924
rect 46987 3896 47032 3924
rect 47026 3884 47032 3896
rect 47084 3884 47090 3936
rect 47578 3884 47584 3936
rect 47636 3924 47642 3936
rect 50154 3924 50160 3936
rect 47636 3896 50160 3924
rect 47636 3884 47642 3896
rect 50154 3884 50160 3896
rect 50212 3884 50218 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2958 3720 2964 3732
rect 2179 3692 2964 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 5261 3723 5319 3729
rect 5261 3689 5273 3723
rect 5307 3720 5319 3723
rect 5350 3720 5356 3732
rect 5307 3692 5356 3720
rect 5307 3689 5319 3692
rect 5261 3683 5319 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 7190 3720 7196 3732
rect 6696 3692 7052 3720
rect 7151 3692 7196 3720
rect 6696 3680 6702 3692
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 6914 3652 6920 3664
rect 6788 3624 6920 3652
rect 6788 3612 6794 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7024 3652 7052 3692
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 9122 3720 9128 3732
rect 7800 3692 9128 3720
rect 7800 3680 7806 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 9416 3692 9505 3720
rect 9416 3664 9444 3692
rect 9493 3689 9505 3692
rect 9539 3689 9551 3723
rect 9493 3683 9551 3689
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 35894 3720 35900 3732
rect 10928 3692 35900 3720
rect 10928 3680 10934 3692
rect 35894 3680 35900 3692
rect 35952 3680 35958 3732
rect 36906 3720 36912 3732
rect 36867 3692 36912 3720
rect 36906 3680 36912 3692
rect 36964 3680 36970 3732
rect 38378 3680 38384 3732
rect 38436 3720 38442 3732
rect 38749 3723 38807 3729
rect 38749 3720 38761 3723
rect 38436 3692 38761 3720
rect 38436 3680 38442 3692
rect 38749 3689 38761 3692
rect 38795 3689 38807 3723
rect 38749 3683 38807 3689
rect 39390 3680 39396 3732
rect 39448 3720 39454 3732
rect 41414 3720 41420 3732
rect 39448 3692 41420 3720
rect 39448 3680 39454 3692
rect 41414 3680 41420 3692
rect 41472 3680 41478 3732
rect 42794 3720 42800 3732
rect 42755 3692 42800 3720
rect 42794 3680 42800 3692
rect 42852 3680 42858 3732
rect 47489 3723 47547 3729
rect 47489 3720 47501 3723
rect 47320 3692 47501 3720
rect 9306 3652 9312 3664
rect 7024 3624 9312 3652
rect 9306 3612 9312 3624
rect 9364 3612 9370 3664
rect 9398 3612 9404 3664
rect 9456 3612 9462 3664
rect 12069 3655 12127 3661
rect 12069 3621 12081 3655
rect 12115 3652 12127 3655
rect 14918 3652 14924 3664
rect 12115 3624 14924 3652
rect 12115 3621 12127 3624
rect 12069 3615 12127 3621
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 16574 3612 16580 3664
rect 16632 3652 16638 3664
rect 16853 3655 16911 3661
rect 16853 3652 16865 3655
rect 16632 3624 16865 3652
rect 16632 3612 16638 3624
rect 16853 3621 16865 3624
rect 16899 3621 16911 3655
rect 20162 3652 20168 3664
rect 16853 3615 16911 3621
rect 17788 3624 20168 3652
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 9214 3584 9220 3596
rect 4479 3556 9220 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 1854 3516 1860 3528
rect 1815 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 2682 3516 2688 3528
rect 2643 3488 2688 3516
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4448 3516 4476 3547
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 12986 3584 12992 3596
rect 12176 3556 12992 3584
rect 3835 3488 4476 3516
rect 4525 3519 4583 3525
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 198 3408 204 3460
rect 256 3448 262 3460
rect 4540 3448 4568 3479
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 5132 3488 5181 3516
rect 5132 3476 5138 3488
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 6641 3519 6699 3525
rect 6641 3516 6653 3519
rect 5592 3488 6653 3516
rect 5592 3476 5598 3488
rect 6641 3485 6653 3488
rect 6687 3516 6699 3519
rect 6730 3516 6736 3528
rect 6687 3488 6736 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 7466 3516 7472 3528
rect 7423 3488 7472 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7834 3516 7840 3528
rect 7795 3488 7840 3516
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8018 3516 8024 3528
rect 7979 3488 8024 3516
rect 8018 3476 8024 3488
rect 8076 3516 8082 3528
rect 8076 3488 9444 3516
rect 8076 3476 8082 3488
rect 9416 3448 9444 3488
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9674 3516 9680 3528
rect 9548 3488 9593 3516
rect 9635 3488 9680 3516
rect 9548 3476 9554 3488
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 10594 3516 10600 3528
rect 9824 3488 9869 3516
rect 10555 3488 10600 3516
rect 9824 3476 9830 3488
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 12176 3516 12204 3556
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 15470 3584 15476 3596
rect 13964 3556 14320 3584
rect 15431 3556 15476 3584
rect 13964 3544 13970 3556
rect 10827 3488 12204 3516
rect 12253 3519 12311 3525
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 12253 3485 12265 3519
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3516 12771 3519
rect 13924 3516 13952 3544
rect 12759 3488 13952 3516
rect 12759 3485 12771 3488
rect 12713 3479 12771 3485
rect 10796 3448 10824 3479
rect 256 3420 2912 3448
rect 4540 3420 9352 3448
rect 9416 3420 10824 3448
rect 256 3408 262 3420
rect 2884 3389 2912 3420
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 3602 3340 3608 3392
rect 3660 3380 3666 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 3660 3352 3985 3380
rect 3660 3340 3666 3352
rect 3973 3349 3985 3352
rect 4019 3349 4031 3383
rect 4614 3380 4620 3392
rect 4575 3352 4620 3380
rect 3973 3343 4031 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 5813 3383 5871 3389
rect 5813 3380 5825 3383
rect 5132 3352 5825 3380
rect 5132 3340 5138 3352
rect 5813 3349 5825 3352
rect 5859 3349 5871 3383
rect 6454 3380 6460 3392
rect 6415 3352 6460 3380
rect 5813 3343 5871 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8662 3380 8668 3392
rect 8251 3352 8668 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 9324 3380 9352 3420
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 10928 3420 11437 3448
rect 10928 3408 10934 3420
rect 11425 3417 11437 3420
rect 11471 3417 11483 3451
rect 12268 3448 12296 3479
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14292 3525 14320 3556
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15746 3525 15752 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 14056 3488 14105 3516
rect 14056 3476 14062 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 15740 3516 15752 3525
rect 15707 3488 15752 3516
rect 14277 3479 14335 3485
rect 15740 3479 15752 3488
rect 15746 3476 15752 3479
rect 15804 3476 15810 3528
rect 17788 3525 17816 3624
rect 20162 3612 20168 3624
rect 20220 3612 20226 3664
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 22094 3652 22100 3664
rect 21876 3624 22100 3652
rect 21876 3612 21882 3624
rect 22094 3612 22100 3624
rect 22152 3612 22158 3664
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 23014 3652 23020 3664
rect 22244 3624 23020 3652
rect 22244 3612 22250 3624
rect 23014 3612 23020 3624
rect 23072 3612 23078 3664
rect 23290 3652 23296 3664
rect 23251 3624 23296 3652
rect 23290 3612 23296 3624
rect 23348 3612 23354 3664
rect 24486 3612 24492 3664
rect 24544 3652 24550 3664
rect 25866 3652 25872 3664
rect 24544 3624 25872 3652
rect 24544 3612 24550 3624
rect 20346 3584 20352 3596
rect 18708 3556 20352 3584
rect 18708 3525 18736 3556
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 24394 3544 24400 3596
rect 24452 3584 24458 3596
rect 25041 3587 25099 3593
rect 24452 3556 24716 3584
rect 24452 3544 24458 3556
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18840 3488 19441 3516
rect 18840 3476 18846 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20254 3476 20260 3528
rect 20312 3516 20318 3528
rect 20441 3519 20499 3525
rect 20441 3516 20453 3519
rect 20312 3488 20453 3516
rect 20312 3476 20318 3488
rect 20441 3485 20453 3488
rect 20487 3516 20499 3519
rect 20530 3516 20536 3528
rect 20487 3488 20536 3516
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 22646 3516 22652 3528
rect 22607 3488 22652 3516
rect 22646 3476 22652 3488
rect 22704 3476 22710 3528
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 23014 3516 23020 3528
rect 22796 3488 22841 3516
rect 22975 3488 23020 3516
rect 22796 3476 22802 3488
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23155 3519 23213 3525
rect 23155 3485 23167 3519
rect 23201 3516 23213 3519
rect 23474 3516 23480 3528
rect 23201 3488 23480 3516
rect 23201 3485 23213 3488
rect 23155 3479 23213 3485
rect 23474 3476 23480 3488
rect 23532 3516 23538 3528
rect 24486 3516 24492 3528
rect 23532 3488 24492 3516
rect 23532 3476 23538 3488
rect 24486 3476 24492 3488
rect 24544 3476 24550 3528
rect 24688 3525 24716 3556
rect 25041 3553 25053 3587
rect 25087 3584 25099 3587
rect 25087 3556 25167 3584
rect 25087 3553 25099 3556
rect 25041 3547 25099 3553
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 24854 3516 24860 3528
rect 24912 3525 24918 3528
rect 24819 3488 24860 3516
rect 24673 3479 24731 3485
rect 24854 3476 24860 3488
rect 24912 3479 24919 3525
rect 24958 3519 25016 3525
rect 24958 3485 24970 3519
rect 25004 3516 25016 3519
rect 25004 3488 25084 3516
rect 25004 3485 25016 3488
rect 24958 3479 25016 3485
rect 24912 3476 24918 3479
rect 13354 3448 13360 3460
rect 12268 3420 13360 3448
rect 11425 3411 11483 3417
rect 13354 3408 13360 3420
rect 13412 3408 13418 3460
rect 17126 3408 17132 3460
rect 17184 3448 17190 3460
rect 20708 3451 20766 3457
rect 17184 3420 20668 3448
rect 17184 3408 17190 3420
rect 10778 3380 10784 3392
rect 9324 3352 10784 3380
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 10962 3380 10968 3392
rect 10923 3352 10968 3380
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 14461 3383 14519 3389
rect 14461 3349 14473 3383
rect 14507 3380 14519 3383
rect 15378 3380 15384 3392
rect 14507 3352 15384 3380
rect 14507 3349 14519 3352
rect 14461 3343 14519 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 17310 3380 17316 3392
rect 15528 3352 17316 3380
rect 15528 3340 15534 3352
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 17678 3340 17684 3392
rect 17736 3380 17742 3392
rect 17957 3383 18015 3389
rect 17957 3380 17969 3383
rect 17736 3352 17969 3380
rect 17736 3340 17742 3352
rect 17957 3349 17969 3352
rect 18003 3349 18015 3383
rect 18506 3380 18512 3392
rect 18467 3352 18512 3380
rect 17957 3343 18015 3349
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 19242 3380 19248 3392
rect 19203 3352 19248 3380
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 20640 3380 20668 3420
rect 20708 3417 20720 3451
rect 20754 3448 20766 3451
rect 21082 3448 21088 3460
rect 20754 3420 21088 3448
rect 20754 3417 20766 3420
rect 20708 3411 20766 3417
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 22922 3448 22928 3460
rect 22883 3420 22928 3448
rect 22922 3408 22928 3420
rect 22980 3408 22986 3460
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 20640 3352 21833 3380
rect 21821 3349 21833 3352
rect 21867 3380 21879 3383
rect 23014 3380 23020 3392
rect 21867 3352 23020 3380
rect 21867 3349 21879 3352
rect 21821 3343 21879 3349
rect 23014 3340 23020 3352
rect 23072 3380 23078 3392
rect 25056 3380 25084 3488
rect 25139 3448 25167 3556
rect 25236 3519 25294 3525
rect 25236 3485 25248 3519
rect 25282 3516 25294 3519
rect 25332 3516 25360 3624
rect 25866 3612 25872 3624
rect 25924 3612 25930 3664
rect 26970 3612 26976 3664
rect 27028 3652 27034 3664
rect 27028 3624 36584 3652
rect 27028 3612 27034 3624
rect 31202 3544 31208 3596
rect 31260 3584 31266 3596
rect 36440 3584 36446 3596
rect 31260 3556 31340 3584
rect 36401 3556 36446 3584
rect 31260 3544 31266 3556
rect 25282 3488 25360 3516
rect 25282 3485 25294 3488
rect 25236 3479 25294 3485
rect 25590 3476 25596 3528
rect 25648 3516 25654 3528
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 25648 3488 25881 3516
rect 25648 3476 25654 3488
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 25869 3479 25927 3485
rect 26136 3519 26194 3525
rect 26136 3485 26148 3519
rect 26182 3516 26194 3519
rect 26418 3516 26424 3528
rect 26182 3488 26424 3516
rect 26182 3485 26194 3488
rect 26136 3479 26194 3485
rect 26418 3476 26424 3488
rect 26476 3476 26482 3528
rect 31021 3519 31079 3525
rect 31021 3485 31033 3519
rect 31067 3516 31079 3519
rect 31110 3516 31116 3528
rect 31067 3488 31116 3516
rect 31067 3485 31079 3488
rect 31021 3479 31079 3485
rect 31110 3476 31116 3488
rect 31168 3476 31174 3528
rect 31312 3525 31340 3556
rect 36440 3544 36446 3556
rect 36498 3544 36504 3596
rect 36556 3584 36584 3624
rect 36722 3612 36728 3664
rect 36780 3652 36786 3664
rect 43438 3652 43444 3664
rect 36780 3624 43444 3652
rect 36780 3612 36786 3624
rect 43438 3612 43444 3624
rect 43496 3612 43502 3664
rect 46382 3612 46388 3664
rect 46440 3652 46446 3664
rect 47320 3652 47348 3692
rect 47489 3689 47501 3692
rect 47535 3689 47547 3723
rect 47489 3683 47547 3689
rect 47578 3680 47584 3732
rect 47636 3720 47642 3732
rect 57146 3720 57152 3732
rect 47636 3692 57152 3720
rect 47636 3680 47642 3692
rect 57146 3680 57152 3692
rect 57204 3680 57210 3732
rect 46440 3624 47348 3652
rect 46440 3612 46446 3624
rect 47946 3612 47952 3664
rect 48004 3652 48010 3664
rect 48004 3624 49096 3652
rect 48004 3612 48010 3624
rect 42150 3584 42156 3596
rect 36556 3556 42156 3584
rect 42150 3544 42156 3556
rect 42208 3544 42214 3596
rect 47578 3544 47584 3596
rect 47636 3584 47642 3596
rect 48498 3584 48504 3596
rect 47636 3556 48504 3584
rect 47636 3544 47642 3556
rect 48498 3544 48504 3556
rect 48556 3544 48562 3596
rect 31297 3519 31355 3525
rect 31297 3485 31309 3519
rect 31343 3485 31355 3519
rect 31297 3479 31355 3485
rect 31389 3519 31447 3525
rect 31389 3485 31401 3519
rect 31435 3516 31447 3519
rect 31570 3516 31576 3528
rect 31435 3488 31576 3516
rect 31435 3485 31447 3488
rect 31389 3479 31447 3485
rect 31570 3476 31576 3488
rect 31628 3476 31634 3528
rect 32122 3516 32128 3528
rect 32083 3488 32128 3516
rect 32122 3476 32128 3488
rect 32180 3476 32186 3528
rect 32232 3488 34744 3516
rect 25774 3448 25780 3460
rect 25139 3420 25780 3448
rect 25774 3408 25780 3420
rect 25832 3408 25838 3460
rect 31202 3448 31208 3460
rect 31163 3420 31208 3448
rect 31202 3408 31208 3420
rect 31260 3408 31266 3460
rect 32232 3448 32260 3488
rect 31404 3420 32260 3448
rect 25406 3380 25412 3392
rect 23072 3352 25084 3380
rect 25367 3352 25412 3380
rect 23072 3340 23078 3352
rect 25406 3340 25412 3352
rect 25464 3340 25470 3392
rect 25958 3340 25964 3392
rect 26016 3380 26022 3392
rect 27249 3383 27307 3389
rect 27249 3380 27261 3383
rect 26016 3352 27261 3380
rect 26016 3340 26022 3352
rect 27249 3349 27261 3352
rect 27295 3349 27307 3383
rect 27249 3343 27307 3349
rect 31110 3340 31116 3392
rect 31168 3380 31174 3392
rect 31404 3380 31432 3420
rect 31570 3380 31576 3392
rect 31168 3352 31432 3380
rect 31531 3352 31576 3380
rect 31168 3340 31174 3352
rect 31570 3340 31576 3352
rect 31628 3340 31634 3392
rect 32232 3389 32260 3420
rect 33505 3451 33563 3457
rect 33505 3417 33517 3451
rect 33551 3448 33563 3451
rect 34422 3448 34428 3460
rect 33551 3420 34428 3448
rect 33551 3417 33563 3420
rect 33505 3411 33563 3417
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 32217 3383 32275 3389
rect 32217 3349 32229 3383
rect 32263 3349 32275 3383
rect 32217 3343 32275 3349
rect 32306 3340 32312 3392
rect 32364 3380 32370 3392
rect 33597 3383 33655 3389
rect 33597 3380 33609 3383
rect 32364 3352 33609 3380
rect 32364 3340 32370 3352
rect 33597 3349 33609 3352
rect 33643 3380 33655 3383
rect 34514 3380 34520 3392
rect 33643 3352 34520 3380
rect 33643 3349 33655 3352
rect 33597 3343 33655 3349
rect 34514 3340 34520 3352
rect 34572 3340 34578 3392
rect 34716 3380 34744 3488
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34848 3488 34897 3516
rect 34848 3476 34854 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 35161 3519 35219 3525
rect 35161 3485 35173 3519
rect 35207 3516 35219 3519
rect 35342 3516 35348 3528
rect 35207 3488 35348 3516
rect 35207 3485 35219 3488
rect 35161 3479 35219 3485
rect 35342 3476 35348 3488
rect 35400 3476 35406 3528
rect 36078 3476 36084 3528
rect 36136 3516 36142 3528
rect 36630 3525 36636 3528
rect 36173 3519 36231 3525
rect 36173 3516 36185 3519
rect 36136 3488 36185 3516
rect 36136 3476 36142 3488
rect 36173 3485 36185 3488
rect 36219 3485 36231 3519
rect 36173 3479 36231 3485
rect 36345 3519 36403 3525
rect 36345 3485 36357 3519
rect 36391 3485 36403 3519
rect 36345 3479 36403 3485
rect 36587 3519 36636 3525
rect 36587 3485 36599 3519
rect 36633 3485 36636 3519
rect 36587 3479 36636 3485
rect 35526 3408 35532 3460
rect 35584 3448 35590 3460
rect 36372 3448 36400 3479
rect 36630 3476 36636 3479
rect 36688 3476 36694 3528
rect 36725 3519 36783 3525
rect 36725 3485 36737 3519
rect 36771 3518 36783 3519
rect 36771 3516 36860 3518
rect 36998 3516 37004 3528
rect 36771 3490 37004 3516
rect 36771 3485 36783 3490
rect 36832 3488 37004 3490
rect 36725 3479 36783 3485
rect 36998 3476 37004 3488
rect 37056 3476 37062 3528
rect 38194 3516 38200 3528
rect 38155 3488 38200 3516
rect 38194 3476 38200 3488
rect 38252 3476 38258 3528
rect 38286 3476 38292 3528
rect 38344 3516 38350 3528
rect 38565 3519 38623 3525
rect 38565 3516 38577 3519
rect 38344 3488 38577 3516
rect 38344 3476 38350 3488
rect 38565 3485 38577 3488
rect 38611 3485 38623 3519
rect 38565 3479 38623 3485
rect 40126 3476 40132 3528
rect 40184 3516 40190 3528
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 40184 3488 40509 3516
rect 40184 3476 40190 3488
rect 40497 3485 40509 3488
rect 40543 3516 40555 3519
rect 40770 3516 40776 3528
rect 40543 3488 40776 3516
rect 40543 3485 40555 3488
rect 40497 3479 40555 3485
rect 40770 3476 40776 3488
rect 40828 3476 40834 3528
rect 41230 3516 41236 3528
rect 41191 3488 41236 3516
rect 41230 3476 41236 3488
rect 41288 3476 41294 3528
rect 41506 3516 41512 3528
rect 41467 3488 41512 3516
rect 41506 3476 41512 3488
rect 41564 3476 41570 3528
rect 41601 3519 41659 3525
rect 41601 3485 41613 3519
rect 41647 3485 41659 3519
rect 42242 3516 42248 3528
rect 42203 3488 42248 3516
rect 41601 3479 41659 3485
rect 38381 3451 38439 3457
rect 38381 3448 38393 3451
rect 35584 3420 36400 3448
rect 36832 3420 38393 3448
rect 35584 3408 35590 3420
rect 36832 3380 36860 3420
rect 38381 3417 38393 3420
rect 38427 3417 38439 3451
rect 38381 3411 38439 3417
rect 38473 3451 38531 3457
rect 38473 3417 38485 3451
rect 38519 3448 38531 3451
rect 39850 3448 39856 3460
rect 38519 3420 39856 3448
rect 38519 3417 38531 3420
rect 38473 3411 38531 3417
rect 34716 3352 36860 3380
rect 38396 3380 38424 3411
rect 39850 3408 39856 3420
rect 39908 3408 39914 3460
rect 41322 3408 41328 3460
rect 41380 3448 41386 3460
rect 41417 3451 41475 3457
rect 41417 3448 41429 3451
rect 41380 3420 41429 3448
rect 41380 3408 41386 3420
rect 41417 3417 41429 3420
rect 41463 3417 41475 3451
rect 41616 3448 41644 3479
rect 42242 3476 42248 3488
rect 42300 3476 42306 3528
rect 42518 3525 42524 3528
rect 42517 3516 42524 3525
rect 42479 3488 42524 3516
rect 42517 3479 42524 3488
rect 42518 3476 42524 3479
rect 42576 3476 42582 3528
rect 42613 3519 42671 3525
rect 42613 3485 42625 3519
rect 42659 3516 42671 3519
rect 42702 3516 42708 3528
rect 42659 3488 42708 3516
rect 42659 3485 42671 3488
rect 42613 3479 42671 3485
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 42794 3476 42800 3528
rect 42852 3516 42858 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 42852 3488 43269 3516
rect 42852 3476 42858 3488
rect 43257 3485 43269 3488
rect 43303 3516 43315 3519
rect 43806 3516 43812 3528
rect 43303 3488 43812 3516
rect 43303 3485 43315 3488
rect 43257 3479 43315 3485
rect 43806 3476 43812 3488
rect 43864 3476 43870 3528
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45922 3516 45928 3528
rect 45883 3488 45928 3516
rect 45922 3476 45928 3488
rect 45980 3476 45986 3528
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3485 46167 3519
rect 46290 3516 46296 3528
rect 46251 3488 46296 3516
rect 46109 3479 46167 3485
rect 41417 3411 41475 3417
rect 41524 3420 41644 3448
rect 42429 3451 42487 3457
rect 39574 3380 39580 3392
rect 38396 3352 39580 3380
rect 39574 3340 39580 3352
rect 39632 3340 39638 3392
rect 39666 3340 39672 3392
rect 39724 3380 39730 3392
rect 40681 3383 40739 3389
rect 40681 3380 40693 3383
rect 39724 3352 40693 3380
rect 39724 3340 39730 3352
rect 40681 3349 40693 3352
rect 40727 3349 40739 3383
rect 40681 3343 40739 3349
rect 40862 3340 40868 3392
rect 40920 3380 40926 3392
rect 41524 3380 41552 3420
rect 42429 3417 42441 3451
rect 42475 3448 42487 3451
rect 46124 3448 46152 3479
rect 46290 3476 46296 3488
rect 46348 3476 46354 3528
rect 46934 3516 46940 3528
rect 46895 3488 46940 3516
rect 46934 3476 46940 3488
rect 46992 3476 46998 3528
rect 47118 3476 47124 3528
rect 47176 3516 47182 3528
rect 47351 3519 47409 3525
rect 47176 3488 47221 3516
rect 47176 3476 47182 3488
rect 47351 3485 47363 3519
rect 47397 3516 47409 3519
rect 47486 3516 47492 3528
rect 47397 3488 47492 3516
rect 47397 3485 47409 3488
rect 47351 3479 47409 3485
rect 47486 3476 47492 3488
rect 47544 3476 47550 3528
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 48866 3516 48872 3528
rect 47912 3488 48872 3516
rect 47912 3476 47918 3488
rect 48866 3476 48872 3488
rect 48924 3476 48930 3528
rect 49068 3525 49096 3624
rect 51166 3544 51172 3596
rect 51224 3584 51230 3596
rect 57977 3587 58035 3593
rect 57977 3584 57989 3587
rect 51224 3556 57989 3584
rect 51224 3544 51230 3556
rect 57977 3553 57989 3556
rect 58023 3553 58035 3587
rect 57977 3547 58035 3553
rect 49053 3519 49111 3525
rect 49053 3485 49065 3519
rect 49099 3485 49111 3519
rect 49053 3479 49111 3485
rect 49252 3488 49433 3516
rect 42475 3420 42564 3448
rect 42475 3417 42487 3420
rect 42429 3411 42487 3417
rect 41782 3380 41788 3392
rect 40920 3352 41552 3380
rect 41743 3352 41788 3380
rect 40920 3340 40926 3352
rect 41782 3340 41788 3352
rect 41840 3340 41846 3392
rect 42536 3380 42564 3420
rect 42812 3420 46152 3448
rect 46201 3451 46259 3457
rect 42702 3380 42708 3392
rect 42536 3352 42708 3380
rect 42702 3340 42708 3352
rect 42760 3380 42766 3392
rect 42812 3380 42840 3420
rect 46201 3417 46213 3451
rect 46247 3448 46259 3451
rect 46658 3448 46664 3460
rect 46247 3420 46664 3448
rect 46247 3417 46259 3420
rect 46201 3411 46259 3417
rect 46658 3408 46664 3420
rect 46716 3408 46722 3460
rect 47210 3408 47216 3460
rect 47268 3448 47274 3460
rect 47268 3420 47313 3448
rect 47268 3408 47274 3420
rect 48038 3408 48044 3460
rect 48096 3448 48102 3460
rect 49252 3448 49280 3488
rect 48096 3420 49280 3448
rect 49405 3448 49433 3488
rect 49602 3476 49608 3528
rect 49660 3516 49666 3528
rect 50157 3519 50215 3525
rect 50157 3516 50169 3519
rect 49660 3488 50169 3516
rect 49660 3476 49666 3488
rect 50157 3485 50169 3488
rect 50203 3485 50215 3519
rect 50157 3479 50215 3485
rect 57701 3519 57759 3525
rect 57701 3485 57713 3519
rect 57747 3516 57759 3519
rect 58158 3516 58164 3528
rect 57747 3488 58164 3516
rect 57747 3485 57759 3488
rect 57701 3479 57759 3485
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 50402 3451 50460 3457
rect 50402 3448 50414 3451
rect 49405 3420 50414 3448
rect 48096 3408 48102 3420
rect 50402 3417 50414 3420
rect 50448 3417 50460 3451
rect 50402 3411 50460 3417
rect 42760 3352 42840 3380
rect 42760 3340 42766 3352
rect 42978 3340 42984 3392
rect 43036 3380 43042 3392
rect 43441 3383 43499 3389
rect 43441 3380 43453 3383
rect 43036 3352 43453 3380
rect 43036 3340 43042 3352
rect 43441 3349 43453 3352
rect 43487 3349 43499 3383
rect 43441 3343 43499 3349
rect 45373 3383 45431 3389
rect 45373 3349 45385 3383
rect 45419 3380 45431 3383
rect 45462 3380 45468 3392
rect 45419 3352 45468 3380
rect 45419 3349 45431 3352
rect 45373 3343 45431 3349
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 46474 3380 46480 3392
rect 46435 3352 46480 3380
rect 46474 3340 46480 3352
rect 46532 3340 46538 3392
rect 46934 3340 46940 3392
rect 46992 3380 46998 3392
rect 48314 3380 48320 3392
rect 46992 3352 48320 3380
rect 46992 3340 46998 3352
rect 48314 3340 48320 3352
rect 48372 3340 48378 3392
rect 48406 3340 48412 3392
rect 48464 3380 48470 3392
rect 49237 3383 49295 3389
rect 49237 3380 49249 3383
rect 48464 3352 49249 3380
rect 48464 3340 48470 3352
rect 49237 3349 49249 3352
rect 49283 3349 49295 3383
rect 51534 3380 51540 3392
rect 51495 3352 51540 3380
rect 49237 3343 49295 3349
rect 51534 3340 51540 3352
rect 51592 3340 51598 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 7285 3179 7343 3185
rect 2179 3148 7236 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 5166 3108 5172 3120
rect 3436 3080 5172 3108
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 3234 3040 3240 3052
rect 2731 3012 3240 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3436 3049 3464 3080
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 6822 3108 6828 3120
rect 6748 3080 6828 3108
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 4700 3043 4758 3049
rect 4700 3009 4712 3043
rect 4746 3040 4758 3043
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 4746 3012 6377 3040
rect 4746 3009 4758 3012
rect 4700 3003 4758 3009
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6365 3003 6423 3009
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6748 3049 6776 3080
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 7208 3108 7236 3148
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 8294 3176 8300 3188
rect 7331 3148 8300 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8444 3148 9536 3176
rect 8444 3136 8450 3148
rect 9398 3117 9404 3120
rect 9392 3108 9404 3117
rect 7208 3080 8800 3108
rect 9359 3080 9404 3108
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6733 3003 6791 3009
rect 7116 3012 7481 3040
rect 1946 2932 1952 2984
rect 2004 2972 2010 2984
rect 3326 2972 3332 2984
rect 2004 2944 3332 2972
rect 2004 2932 2010 2944
rect 3326 2932 3332 2944
rect 3384 2972 3390 2984
rect 3786 2972 3792 2984
rect 3384 2944 3792 2972
rect 3384 2932 3390 2944
rect 3786 2932 3792 2944
rect 3844 2972 3850 2984
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 3844 2944 4445 2972
rect 3844 2932 3850 2944
rect 4433 2941 4445 2944
rect 4479 2941 4491 2975
rect 4433 2935 4491 2941
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5500 2944 6837 2972
rect 5500 2932 5506 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 716 2876 3617 2904
rect 716 2864 722 2876
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 7116 2904 7144 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 8386 3040 8392 3052
rect 7616 3012 8392 3040
rect 7616 3000 7622 3012
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 8772 3040 8800 3080
rect 9392 3071 9404 3080
rect 9398 3068 9404 3071
rect 9456 3068 9462 3120
rect 9508 3108 9536 3148
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 9640 3148 10517 3176
rect 9640 3136 9646 3148
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 10505 3139 10563 3145
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 15102 3176 15108 3188
rect 14139 3148 15108 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15841 3179 15899 3185
rect 15841 3145 15853 3179
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 12897 3111 12955 3117
rect 9508 3080 12434 3108
rect 9950 3040 9956 3052
rect 8772 3012 9956 3040
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11020 3012 11713 3040
rect 11020 3000 11026 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 12406 3040 12434 3080
rect 12897 3077 12909 3111
rect 12943 3108 12955 3111
rect 12943 3080 14780 3108
rect 12943 3077 12955 3080
rect 12897 3071 12955 3077
rect 12529 3043 12587 3049
rect 12529 3040 12541 3043
rect 12406 3012 12541 3040
rect 11701 3003 11759 3009
rect 12529 3009 12541 3012
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12986 3040 12992 3052
rect 12759 3012 12992 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14752 3049 14780 3080
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 14737 3003 14795 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8312 2944 9137 2972
rect 3605 2867 3663 2873
rect 5368 2876 7144 2904
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 2648 2808 2881 2836
rect 2648 2796 2654 2808
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 2869 2799 2927 2805
rect 4706 2796 4712 2848
rect 4764 2836 4770 2848
rect 5368 2836 5396 2876
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 8312 2904 8340 2944
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 13725 2975 13783 2981
rect 10192 2944 12434 2972
rect 10192 2932 10198 2944
rect 7340 2876 8340 2904
rect 12406 2904 12434 2944
rect 13725 2941 13737 2975
rect 13771 2941 13783 2975
rect 15856 2972 15884 3139
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 19392 3148 19717 3176
rect 19392 3136 19398 3148
rect 19705 3145 19717 3148
rect 19751 3176 19763 3179
rect 19978 3176 19984 3188
rect 19751 3148 19984 3176
rect 19751 3145 19763 3148
rect 19705 3139 19763 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 20070 3136 20076 3188
rect 20128 3176 20134 3188
rect 20441 3179 20499 3185
rect 20441 3176 20453 3179
rect 20128 3148 20453 3176
rect 20128 3136 20134 3148
rect 20441 3145 20453 3148
rect 20487 3145 20499 3179
rect 21082 3176 21088 3188
rect 21043 3148 21088 3176
rect 20441 3139 20499 3145
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 22370 3136 22376 3188
rect 22428 3176 22434 3188
rect 24854 3176 24860 3188
rect 22428 3148 24860 3176
rect 22428 3136 22434 3148
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 25590 3176 25596 3188
rect 25056 3148 25596 3176
rect 17310 3068 17316 3120
rect 17368 3108 17374 3120
rect 18592 3111 18650 3117
rect 17368 3080 18092 3108
rect 17368 3068 17374 3080
rect 16022 3040 16028 3052
rect 15983 3012 16028 3040
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17494 3040 17500 3052
rect 16899 3012 17500 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 17604 2972 17632 3003
rect 15856 2944 17632 2972
rect 18064 2972 18092 3080
rect 18592 3077 18604 3111
rect 18638 3108 18650 3111
rect 18966 3108 18972 3120
rect 18638 3080 18972 3108
rect 18638 3077 18650 3080
rect 18592 3071 18650 3077
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 22002 3068 22008 3120
rect 22060 3108 22066 3120
rect 23014 3108 23020 3120
rect 22060 3080 22784 3108
rect 22975 3080 23020 3108
rect 22060 3068 22066 3080
rect 20254 3040 20260 3052
rect 18432 3012 20260 3040
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 18064 2944 18337 2972
rect 13725 2935 13783 2941
rect 18325 2941 18337 2944
rect 18371 2972 18383 2975
rect 18432 2972 18460 3012
rect 20254 3000 20260 3012
rect 20312 3000 20318 3052
rect 20625 3043 20683 3049
rect 20625 3009 20637 3043
rect 20671 3040 20683 3043
rect 21082 3040 21088 3052
rect 20671 3012 21088 3040
rect 20671 3009 20683 3012
rect 20625 3003 20683 3009
rect 21082 3000 21088 3012
rect 21140 3000 21146 3052
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21818 3040 21824 3052
rect 21779 3012 21824 3040
rect 21269 3003 21327 3009
rect 18371 2944 18460 2972
rect 21284 2972 21312 3003
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22646 3040 22652 3052
rect 22607 3012 22652 3040
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 22756 3049 22784 3080
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 25056 3108 25084 3148
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 25682 3136 25688 3188
rect 25740 3176 25746 3188
rect 26973 3179 27031 3185
rect 26973 3176 26985 3179
rect 25740 3148 26985 3176
rect 25740 3136 25746 3148
rect 26973 3145 26985 3148
rect 27019 3145 27031 3179
rect 26973 3139 27031 3145
rect 27246 3136 27252 3188
rect 27304 3176 27310 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 27304 3148 27629 3176
rect 27304 3136 27310 3148
rect 27617 3145 27629 3148
rect 27663 3145 27675 3179
rect 31018 3176 31024 3188
rect 27617 3139 27675 3145
rect 27724 3148 31024 3176
rect 24872 3080 25084 3108
rect 25124 3111 25182 3117
rect 22742 3043 22800 3049
rect 22742 3009 22754 3043
rect 22788 3009 22800 3043
rect 22922 3040 22928 3052
rect 22883 3012 22928 3040
rect 22742 3003 22800 3009
rect 22922 3000 22928 3012
rect 22980 3000 22986 3052
rect 23155 3043 23213 3049
rect 23155 3009 23167 3043
rect 23201 3040 23213 3043
rect 23474 3040 23480 3052
rect 23201 3012 23480 3040
rect 23201 3009 23213 3012
rect 23155 3003 23213 3009
rect 23474 3000 23480 3012
rect 23532 3000 23538 3052
rect 23750 3040 23756 3052
rect 23711 3012 23756 3040
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24118 3000 24124 3052
rect 24176 3040 24182 3052
rect 24872 3049 24900 3080
rect 25124 3077 25136 3111
rect 25170 3108 25182 3111
rect 25406 3108 25412 3120
rect 25170 3080 25412 3108
rect 25170 3077 25182 3080
rect 25124 3071 25182 3077
rect 25406 3068 25412 3080
rect 25464 3068 25470 3120
rect 27724 3108 27752 3148
rect 31018 3136 31024 3148
rect 31076 3136 31082 3188
rect 31202 3136 31208 3188
rect 31260 3176 31266 3188
rect 31481 3179 31539 3185
rect 31481 3176 31493 3179
rect 31260 3148 31493 3176
rect 31260 3136 31266 3148
rect 31481 3145 31493 3148
rect 31527 3145 31539 3179
rect 31481 3139 31539 3145
rect 31846 3136 31852 3188
rect 31904 3176 31910 3188
rect 31904 3148 34008 3176
rect 31904 3136 31910 3148
rect 25516 3080 27752 3108
rect 29356 3111 29414 3117
rect 24857 3043 24915 3049
rect 24857 3040 24869 3043
rect 24176 3012 24869 3040
rect 24176 3000 24182 3012
rect 24857 3009 24869 3012
rect 24903 3009 24915 3043
rect 25516 3040 25544 3080
rect 29356 3077 29368 3111
rect 29402 3108 29414 3111
rect 31386 3108 31392 3120
rect 29402 3080 31392 3108
rect 29402 3077 29414 3080
rect 29356 3071 29414 3077
rect 31386 3068 31392 3080
rect 31444 3068 31450 3120
rect 33680 3111 33738 3117
rect 33680 3077 33692 3111
rect 33726 3108 33738 3111
rect 33870 3108 33876 3120
rect 33726 3080 33876 3108
rect 33726 3077 33738 3080
rect 33680 3071 33738 3077
rect 33870 3068 33876 3080
rect 33928 3068 33934 3120
rect 33980 3108 34008 3148
rect 34698 3136 34704 3188
rect 34756 3176 34762 3188
rect 34793 3179 34851 3185
rect 34793 3176 34805 3179
rect 34756 3148 34805 3176
rect 34756 3136 34762 3148
rect 34793 3145 34805 3148
rect 34839 3145 34851 3179
rect 39390 3176 39396 3188
rect 34793 3139 34851 3145
rect 34900 3148 39396 3176
rect 34900 3108 34928 3148
rect 39390 3136 39396 3148
rect 39448 3136 39454 3188
rect 39577 3179 39635 3185
rect 39577 3145 39589 3179
rect 39623 3176 39635 3179
rect 39850 3176 39856 3188
rect 39623 3148 39856 3176
rect 39623 3145 39635 3148
rect 39577 3139 39635 3145
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 41322 3176 41328 3188
rect 41283 3148 41328 3176
rect 41322 3136 41328 3148
rect 41380 3136 41386 3188
rect 42242 3176 42248 3188
rect 41708 3148 42248 3176
rect 33980 3080 34928 3108
rect 35520 3111 35578 3117
rect 35520 3077 35532 3111
rect 35566 3108 35578 3111
rect 36906 3108 36912 3120
rect 35566 3080 36912 3108
rect 35566 3077 35578 3080
rect 35520 3071 35578 3077
rect 36906 3068 36912 3080
rect 36964 3068 36970 3120
rect 38464 3111 38522 3117
rect 37016 3080 38332 3108
rect 24857 3003 24915 3009
rect 24964 3012 25544 3040
rect 22462 2972 22468 2984
rect 21284 2944 22468 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 13740 2904 13768 2935
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 24964 2972 24992 3012
rect 25958 3000 25964 3052
rect 26016 3040 26022 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26016 3012 27169 3040
rect 26016 3000 26022 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27430 3000 27436 3052
rect 27488 3040 27494 3052
rect 27801 3043 27859 3049
rect 27801 3040 27813 3043
rect 27488 3012 27813 3040
rect 27488 3000 27494 3012
rect 27801 3009 27813 3012
rect 27847 3009 27859 3043
rect 29086 3040 29092 3052
rect 29047 3012 29092 3040
rect 27801 3003 27859 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 30834 3000 30840 3052
rect 30892 3040 30898 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30892 3012 30941 3040
rect 30892 3000 30898 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 31110 3040 31116 3052
rect 31071 3012 31116 3040
rect 30929 3003 30987 3009
rect 31110 3000 31116 3012
rect 31168 3000 31174 3052
rect 31205 3043 31263 3049
rect 31205 3009 31217 3043
rect 31251 3009 31263 3043
rect 31205 3003 31263 3009
rect 31297 3043 31355 3049
rect 31297 3009 31309 3043
rect 31343 3040 31355 3043
rect 32398 3040 32404 3052
rect 31343 3012 31524 3040
rect 32359 3012 32404 3040
rect 31343 3009 31355 3012
rect 31297 3003 31355 3009
rect 22572 2944 24992 2972
rect 12406 2876 13768 2904
rect 7340 2864 7346 2876
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 22572 2904 22600 2944
rect 30282 2932 30288 2984
rect 30340 2972 30346 2984
rect 31220 2972 31248 3003
rect 30340 2944 31248 2972
rect 31496 2972 31524 3012
rect 32398 3000 32404 3012
rect 32456 3000 32462 3052
rect 33410 3040 33416 3052
rect 33323 3012 33416 3040
rect 33410 3000 33416 3012
rect 33468 3040 33474 3052
rect 33468 3012 34468 3040
rect 33468 3000 33474 3012
rect 31938 2972 31944 2984
rect 31496 2944 31944 2972
rect 30340 2932 30346 2944
rect 31938 2932 31944 2944
rect 31996 2972 32002 2984
rect 32306 2972 32312 2984
rect 31996 2944 32312 2972
rect 31996 2932 32002 2944
rect 32306 2932 32312 2944
rect 32364 2932 32370 2984
rect 34440 2972 34468 3012
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 37016 3040 37044 3080
rect 38304 3052 38332 3080
rect 38464 3077 38476 3111
rect 38510 3108 38522 3111
rect 38838 3108 38844 3120
rect 38510 3080 38844 3108
rect 38510 3077 38522 3080
rect 38464 3071 38522 3077
rect 38838 3068 38844 3080
rect 38896 3068 38902 3120
rect 41046 3068 41052 3120
rect 41104 3108 41110 3120
rect 41708 3108 41736 3148
rect 42242 3136 42248 3148
rect 42300 3176 42306 3188
rect 43809 3179 43867 3185
rect 43809 3176 43821 3179
rect 42300 3148 43821 3176
rect 42300 3136 42306 3148
rect 43809 3145 43821 3148
rect 43855 3145 43867 3179
rect 43809 3139 43867 3145
rect 48682 3136 48688 3188
rect 48740 3176 48746 3188
rect 50525 3179 50583 3185
rect 50525 3176 50537 3179
rect 48740 3148 50537 3176
rect 48740 3136 48746 3148
rect 50525 3145 50537 3148
rect 50571 3176 50583 3179
rect 59630 3176 59636 3188
rect 50571 3148 51764 3176
rect 50571 3145 50583 3148
rect 50525 3139 50583 3145
rect 41104 3080 41736 3108
rect 41104 3068 41110 3080
rect 41782 3068 41788 3120
rect 41840 3108 41846 3120
rect 42674 3111 42732 3117
rect 42674 3108 42686 3111
rect 41840 3080 42686 3108
rect 41840 3068 41846 3080
rect 42674 3077 42686 3080
rect 42720 3077 42732 3111
rect 42674 3071 42732 3077
rect 47026 3068 47032 3120
rect 47084 3108 47090 3120
rect 49390 3111 49448 3117
rect 49390 3108 49402 3111
rect 47084 3080 49402 3108
rect 47084 3068 47090 3080
rect 49390 3077 49402 3080
rect 49436 3077 49448 3111
rect 49390 3071 49448 3077
rect 49602 3068 49608 3120
rect 49660 3068 49666 3120
rect 34572 3012 37044 3040
rect 37277 3043 37335 3049
rect 34572 3000 34578 3012
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 38102 3040 38108 3052
rect 37323 3012 38108 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 38102 3000 38108 3012
rect 38160 3000 38166 3052
rect 38286 3000 38292 3052
rect 38344 3040 38350 3052
rect 38344 3012 39804 3040
rect 38344 3000 38350 3012
rect 35250 2972 35256 2984
rect 34440 2944 35256 2972
rect 35250 2932 35256 2944
rect 35308 2932 35314 2984
rect 37918 2932 37924 2984
rect 37976 2972 37982 2984
rect 38197 2975 38255 2981
rect 38197 2972 38209 2975
rect 37976 2944 38209 2972
rect 37976 2932 37982 2944
rect 38197 2941 38209 2944
rect 38243 2941 38255 2975
rect 39776 2972 39804 3012
rect 39850 3000 39856 3052
rect 39908 3040 39914 3052
rect 40037 3043 40095 3049
rect 40037 3040 40049 3043
rect 39908 3012 40049 3040
rect 39908 3000 39914 3012
rect 40037 3009 40049 3012
rect 40083 3009 40095 3043
rect 40770 3040 40776 3052
rect 40731 3012 40776 3040
rect 40037 3003 40095 3009
rect 40770 3000 40776 3012
rect 40828 3000 40834 3052
rect 40862 3000 40868 3052
rect 40920 3040 40926 3052
rect 40957 3043 41015 3049
rect 40957 3040 40969 3043
rect 40920 3012 40969 3040
rect 40920 3000 40926 3012
rect 40957 3009 40969 3012
rect 41003 3009 41015 3043
rect 40957 3003 41015 3009
rect 41138 3000 41144 3052
rect 41196 3040 41202 3052
rect 41196 3012 41241 3040
rect 41196 3000 41202 3012
rect 43898 3000 43904 3052
rect 43956 3040 43962 3052
rect 44269 3043 44327 3049
rect 44269 3040 44281 3043
rect 43956 3012 44281 3040
rect 43956 3000 43962 3012
rect 44269 3009 44281 3012
rect 44315 3009 44327 3043
rect 45646 3040 45652 3052
rect 45607 3012 45652 3040
rect 44269 3003 44327 3009
rect 45646 3000 45652 3012
rect 45704 3000 45710 3052
rect 45922 3049 45928 3052
rect 45916 3003 45928 3049
rect 45980 3040 45986 3052
rect 47581 3043 47639 3049
rect 45980 3012 46016 3040
rect 45922 3000 45928 3003
rect 45980 3000 45986 3012
rect 47581 3009 47593 3043
rect 47627 3040 47639 3043
rect 47762 3040 47768 3052
rect 47627 3012 47768 3040
rect 47627 3009 47639 3012
rect 47581 3003 47639 3009
rect 47762 3000 47768 3012
rect 47820 3000 47826 3052
rect 48590 3000 48596 3052
rect 48648 3040 48654 3052
rect 49145 3043 49203 3049
rect 49145 3040 49157 3043
rect 48648 3012 49157 3040
rect 48648 3000 48654 3012
rect 49145 3009 49157 3012
rect 49191 3040 49203 3043
rect 49620 3040 49648 3068
rect 49191 3012 49648 3040
rect 49191 3009 49203 3012
rect 49145 3003 49203 3009
rect 50154 3000 50160 3052
rect 50212 3040 50218 3052
rect 51736 3049 51764 3148
rect 56888 3148 59636 3176
rect 50985 3043 51043 3049
rect 50985 3040 50997 3043
rect 50212 3012 50997 3040
rect 50212 3000 50218 3012
rect 50985 3009 50997 3012
rect 51031 3009 51043 3043
rect 50985 3003 51043 3009
rect 51721 3043 51779 3049
rect 51721 3009 51733 3043
rect 51767 3009 51779 3043
rect 51721 3003 51779 3009
rect 52178 3000 52184 3052
rect 52236 3040 52242 3052
rect 52917 3043 52975 3049
rect 52917 3040 52929 3043
rect 52236 3012 52929 3040
rect 52236 3000 52242 3012
rect 52917 3009 52929 3012
rect 52963 3009 52975 3043
rect 52917 3003 52975 3009
rect 54389 3043 54447 3049
rect 54389 3009 54401 3043
rect 54435 3009 54447 3043
rect 55858 3040 55864 3052
rect 55819 3012 55864 3040
rect 54389 3003 54447 3009
rect 42426 2972 42432 2984
rect 39776 2944 40908 2972
rect 42387 2944 42432 2972
rect 38197 2935 38255 2941
rect 14884 2876 17908 2904
rect 14884 2864 14890 2876
rect 4764 2808 5396 2836
rect 4764 2796 4770 2808
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5813 2839 5871 2845
rect 5813 2836 5825 2839
rect 5500 2808 5825 2836
rect 5500 2796 5506 2808
rect 5813 2805 5825 2808
rect 5859 2805 5871 2839
rect 5813 2799 5871 2805
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 9766 2836 9772 2848
rect 8527 2808 9772 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12250 2836 12256 2848
rect 11563 2808 12256 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 14553 2839 14611 2845
rect 14553 2805 14565 2839
rect 14599 2836 14611 2839
rect 15102 2836 15108 2848
rect 14599 2808 15108 2836
rect 14599 2805 14611 2808
rect 14553 2799 14611 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15252 2808 15297 2836
rect 15252 2796 15258 2808
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16816 2808 17049 2836
rect 16816 2796 16822 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 17276 2808 17785 2836
rect 17276 2796 17282 2808
rect 17773 2805 17785 2808
rect 17819 2805 17831 2839
rect 17880 2836 17908 2876
rect 19260 2876 22600 2904
rect 19260 2836 19288 2876
rect 22646 2864 22652 2916
rect 22704 2904 22710 2916
rect 23937 2907 23995 2913
rect 23937 2904 23949 2907
rect 22704 2876 23949 2904
rect 22704 2864 22710 2876
rect 23937 2873 23949 2876
rect 23983 2873 23995 2907
rect 36998 2904 37004 2916
rect 23937 2867 23995 2873
rect 25792 2876 26372 2904
rect 17880 2808 19288 2836
rect 17773 2799 17831 2805
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21692 2808 22017 2836
rect 21692 2796 21698 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22922 2796 22928 2848
rect 22980 2836 22986 2848
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 22980 2808 23305 2836
rect 22980 2796 22986 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 23750 2796 23756 2848
rect 23808 2836 23814 2848
rect 25130 2836 25136 2848
rect 23808 2808 25136 2836
rect 23808 2796 23814 2808
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 25590 2796 25596 2848
rect 25648 2836 25654 2848
rect 25792 2836 25820 2876
rect 25648 2808 25820 2836
rect 25648 2796 25654 2808
rect 25866 2796 25872 2848
rect 25924 2836 25930 2848
rect 26237 2839 26295 2845
rect 26237 2836 26249 2839
rect 25924 2808 26249 2836
rect 25924 2796 25930 2808
rect 26237 2805 26249 2808
rect 26283 2805 26295 2839
rect 26344 2836 26372 2876
rect 30208 2876 33456 2904
rect 30208 2836 30236 2876
rect 26344 2808 30236 2836
rect 26237 2799 26295 2805
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30469 2839 30527 2845
rect 30469 2836 30481 2839
rect 30340 2808 30481 2836
rect 30340 2796 30346 2808
rect 30469 2805 30481 2808
rect 30515 2805 30527 2839
rect 30469 2799 30527 2805
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 32585 2839 32643 2845
rect 32585 2836 32597 2839
rect 32364 2808 32597 2836
rect 32364 2796 32370 2808
rect 32585 2805 32597 2808
rect 32631 2805 32643 2839
rect 33428 2836 33456 2876
rect 36648 2876 37004 2904
rect 36648 2845 36676 2876
rect 36998 2864 37004 2876
rect 37056 2864 37062 2916
rect 40221 2907 40279 2913
rect 40221 2904 40233 2907
rect 39132 2876 40233 2904
rect 36633 2839 36691 2845
rect 36633 2836 36645 2839
rect 33428 2808 36645 2836
rect 32585 2799 32643 2805
rect 36633 2805 36645 2808
rect 36679 2805 36691 2839
rect 36633 2799 36691 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36780 2808 37473 2836
rect 36780 2796 36786 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 38194 2796 38200 2848
rect 38252 2836 38258 2848
rect 39132 2836 39160 2876
rect 40221 2873 40233 2876
rect 40267 2873 40279 2907
rect 40880 2904 40908 2944
rect 42426 2932 42432 2944
rect 42484 2932 42490 2984
rect 46750 2932 46756 2984
rect 46808 2972 46814 2984
rect 46808 2944 48912 2972
rect 46808 2932 46814 2944
rect 41138 2904 41144 2916
rect 40880 2876 41144 2904
rect 40221 2867 40279 2873
rect 41138 2864 41144 2876
rect 41196 2864 41202 2916
rect 46934 2864 46940 2916
rect 46992 2904 46998 2916
rect 47765 2907 47823 2913
rect 47765 2904 47777 2907
rect 46992 2876 47777 2904
rect 46992 2864 46998 2876
rect 47765 2873 47777 2876
rect 47811 2873 47823 2907
rect 47765 2867 47823 2873
rect 38252 2808 39160 2836
rect 41156 2836 41184 2864
rect 42610 2836 42616 2848
rect 41156 2808 42616 2836
rect 38252 2796 38258 2808
rect 42610 2796 42616 2808
rect 42668 2796 42674 2848
rect 44082 2796 44088 2848
rect 44140 2836 44146 2848
rect 44453 2839 44511 2845
rect 44453 2836 44465 2839
rect 44140 2808 44465 2836
rect 44140 2796 44146 2808
rect 44453 2805 44465 2808
rect 44499 2805 44511 2839
rect 44453 2799 44511 2805
rect 45646 2796 45652 2848
rect 45704 2836 45710 2848
rect 46382 2836 46388 2848
rect 45704 2808 46388 2836
rect 45704 2796 45710 2808
rect 46382 2796 46388 2808
rect 46440 2796 46446 2848
rect 46658 2796 46664 2848
rect 46716 2836 46722 2848
rect 47029 2839 47087 2845
rect 47029 2836 47041 2839
rect 46716 2808 47041 2836
rect 46716 2796 46722 2808
rect 47029 2805 47041 2808
rect 47075 2836 47087 2839
rect 48774 2836 48780 2848
rect 47075 2808 48780 2836
rect 47075 2805 47087 2808
rect 47029 2799 47087 2805
rect 48774 2796 48780 2808
rect 48832 2796 48838 2848
rect 48884 2836 48912 2944
rect 51534 2932 51540 2984
rect 51592 2972 51598 2984
rect 54404 2972 54432 3003
rect 55858 3000 55864 3012
rect 55916 3000 55922 3052
rect 56888 3049 56916 3148
rect 59630 3136 59636 3148
rect 59688 3136 59694 3188
rect 57146 3108 57152 3120
rect 57107 3080 57152 3108
rect 57146 3068 57152 3080
rect 57204 3068 57210 3120
rect 56873 3043 56931 3049
rect 56873 3009 56885 3043
rect 56919 3009 56931 3043
rect 57885 3043 57943 3049
rect 57885 3040 57897 3043
rect 56873 3003 56931 3009
rect 56980 3012 57897 3040
rect 56980 2972 57008 3012
rect 57885 3009 57897 3012
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 51592 2944 54432 2972
rect 55186 2944 57008 2972
rect 51592 2932 51598 2944
rect 50154 2864 50160 2916
rect 50212 2904 50218 2916
rect 51169 2907 51227 2913
rect 51169 2904 51181 2907
rect 50212 2876 51181 2904
rect 50212 2864 50218 2876
rect 51169 2873 51181 2876
rect 51215 2873 51227 2907
rect 55186 2904 55214 2944
rect 51169 2867 51227 2873
rect 51276 2876 55214 2904
rect 51276 2836 51304 2876
rect 48884 2808 51304 2836
rect 51350 2796 51356 2848
rect 51408 2836 51414 2848
rect 51905 2839 51963 2845
rect 51905 2836 51917 2839
rect 51408 2808 51917 2836
rect 51408 2796 51414 2808
rect 51905 2805 51917 2808
rect 51951 2805 51963 2839
rect 51905 2799 51963 2805
rect 52822 2796 52828 2848
rect 52880 2836 52886 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 52880 2808 53113 2836
rect 52880 2796 52886 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 54294 2796 54300 2848
rect 54352 2836 54358 2848
rect 54573 2839 54631 2845
rect 54573 2836 54585 2839
rect 54352 2808 54585 2836
rect 54352 2796 54358 2808
rect 54573 2805 54585 2808
rect 54619 2805 54631 2839
rect 54573 2799 54631 2805
rect 55766 2796 55772 2848
rect 55824 2836 55830 2848
rect 56045 2839 56103 2845
rect 56045 2836 56057 2839
rect 55824 2808 56057 2836
rect 55824 2796 55830 2808
rect 56045 2805 56057 2808
rect 56091 2805 56103 2839
rect 56045 2799 56103 2805
rect 58069 2839 58127 2845
rect 58069 2805 58081 2839
rect 58115 2836 58127 2839
rect 58710 2836 58716 2848
rect 58115 2808 58716 2836
rect 58115 2805 58127 2808
rect 58069 2799 58127 2805
rect 58710 2796 58716 2808
rect 58768 2796 58774 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 3694 2592 3700 2644
rect 3752 2632 3758 2644
rect 4890 2632 4896 2644
rect 3752 2604 4896 2632
rect 3752 2592 3758 2604
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 11882 2632 11888 2644
rect 8956 2604 11888 2632
rect 1118 2524 1124 2576
rect 1176 2564 1182 2576
rect 4709 2567 4767 2573
rect 4709 2564 4721 2567
rect 1176 2536 4721 2564
rect 1176 2524 1182 2536
rect 4709 2533 4721 2536
rect 4755 2533 4767 2567
rect 4709 2527 4767 2533
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 6549 2567 6607 2573
rect 6549 2564 6561 2567
rect 5592 2536 6561 2564
rect 5592 2524 5598 2536
rect 6549 2533 6561 2536
rect 6595 2533 6607 2567
rect 6549 2527 6607 2533
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3326 2496 3332 2508
rect 3283 2468 3332 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 6270 2496 6276 2508
rect 3804 2468 6276 2496
rect 3804 2437 3832 2468
rect 6270 2456 6276 2468
rect 6328 2456 6334 2508
rect 8846 2496 8852 2508
rect 6380 2468 8852 2496
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4614 2428 4620 2440
rect 4571 2400 4620 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 6380 2437 6408 2468
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 7098 2428 7104 2440
rect 7059 2400 7104 2428
rect 6365 2391 6423 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 1360 2332 1501 2360
rect 1360 2320 1366 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 5552 2360 5580 2391
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 8956 2437 8984 2604
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 19334 2632 19340 2644
rect 14292 2604 19340 2632
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 10597 2567 10655 2573
rect 10597 2564 10609 2567
rect 9456 2536 10609 2564
rect 9456 2524 9462 2536
rect 10597 2533 10609 2536
rect 10643 2533 10655 2567
rect 10597 2527 10655 2533
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 12400 2536 13185 2564
rect 12400 2524 12406 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 13173 2527 13231 2533
rect 14292 2496 14320 2604
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 22186 2632 22192 2644
rect 19444 2604 22192 2632
rect 19444 2564 19472 2604
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 22462 2592 22468 2644
rect 22520 2632 22526 2644
rect 22741 2635 22799 2641
rect 22741 2632 22753 2635
rect 22520 2604 22753 2632
rect 22520 2592 22526 2604
rect 22741 2601 22753 2604
rect 22787 2601 22799 2635
rect 22741 2595 22799 2601
rect 22830 2592 22836 2644
rect 22888 2632 22894 2644
rect 25590 2632 25596 2644
rect 22888 2604 25596 2632
rect 22888 2592 22894 2604
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 28813 2635 28871 2641
rect 28813 2601 28825 2635
rect 28859 2632 28871 2635
rect 28902 2632 28908 2644
rect 28859 2604 28908 2632
rect 28859 2601 28871 2604
rect 28813 2595 28871 2601
rect 28902 2592 28908 2604
rect 28960 2592 28966 2644
rect 30098 2592 30104 2644
rect 30156 2632 30162 2644
rect 30285 2635 30343 2641
rect 30285 2632 30297 2635
rect 30156 2604 30297 2632
rect 30156 2592 30162 2604
rect 30285 2601 30297 2604
rect 30331 2601 30343 2635
rect 30285 2595 30343 2601
rect 34606 2592 34612 2644
rect 34664 2632 34670 2644
rect 34664 2604 35112 2632
rect 34664 2592 34670 2604
rect 18616 2536 19472 2564
rect 15286 2496 15292 2508
rect 11532 2468 14320 2496
rect 14384 2468 15292 2496
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9766 2428 9772 2440
rect 9723 2400 9772 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 11532 2437 11560 2468
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 12250 2428 12256 2440
rect 12211 2400 12256 2428
rect 11517 2391 11575 2397
rect 8754 2360 8760 2372
rect 5552 2332 8760 2360
rect 1489 2323 1547 2329
rect 8754 2320 8760 2332
rect 8812 2320 8818 2372
rect 10428 2360 10456 2391
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 14384 2437 14412 2468
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 15102 2428 15108 2440
rect 15063 2400 15108 2428
rect 14369 2391 14427 2397
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 17126 2428 17132 2440
rect 15887 2400 17132 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17310 2428 17316 2440
rect 17267 2400 17316 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 17488 2431 17546 2437
rect 17488 2397 17500 2431
rect 17534 2428 17546 2431
rect 18506 2428 18512 2440
rect 17534 2400 18512 2428
rect 17534 2397 17546 2400
rect 17488 2391 17546 2397
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 18616 2360 18644 2536
rect 22094 2524 22100 2576
rect 22152 2564 22158 2576
rect 23385 2567 23443 2573
rect 23385 2564 23397 2567
rect 22152 2536 23397 2564
rect 22152 2524 22158 2536
rect 23385 2533 23397 2536
rect 23431 2533 23443 2567
rect 23385 2527 23443 2533
rect 25038 2524 25044 2576
rect 25096 2564 25102 2576
rect 26053 2567 26111 2573
rect 26053 2564 26065 2567
rect 25096 2536 26065 2564
rect 25096 2524 25102 2536
rect 26053 2533 26065 2536
rect 26099 2533 26111 2567
rect 30834 2564 30840 2576
rect 26053 2527 26111 2533
rect 26988 2536 30840 2564
rect 20898 2496 20904 2508
rect 19260 2468 20904 2496
rect 19260 2437 19288 2468
rect 20898 2456 20904 2468
rect 20956 2456 20962 2508
rect 22370 2496 22376 2508
rect 22331 2468 22376 2496
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 22557 2431 22615 2437
rect 20763 2400 22094 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 10428 2332 18644 2360
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3108 2264 3985 2292
rect 3108 2252 3114 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 5721 2295 5779 2301
rect 5721 2261 5733 2295
rect 5767 2292 5779 2295
rect 5994 2292 6000 2304
rect 5767 2264 6000 2292
rect 5767 2261 5779 2264
rect 5721 2255 5779 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 6788 2264 7297 2292
rect 6788 2252 6794 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7984 2264 8033 2292
rect 7984 2252 7990 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8478 2252 8484 2304
rect 8536 2292 8542 2304
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8536 2264 9137 2292
rect 8536 2252 8542 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9272 2264 9873 2292
rect 9272 2252 9278 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 11330 2252 11336 2304
rect 11388 2292 11394 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 11388 2264 11713 2292
rect 11388 2252 11394 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 11940 2264 12449 2292
rect 11940 2252 11946 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 14553 2295 14611 2301
rect 14553 2292 14565 2295
rect 14332 2264 14565 2292
rect 14332 2252 14338 2264
rect 14553 2261 14565 2264
rect 14599 2261 14611 2295
rect 14553 2255 14611 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 14884 2264 15301 2292
rect 14884 2252 14890 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 18616 2301 18644 2332
rect 19058 2320 19064 2372
rect 19116 2360 19122 2372
rect 19996 2360 20024 2391
rect 19116 2332 20024 2360
rect 22066 2360 22094 2400
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 22922 2428 22928 2440
rect 22603 2400 22928 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 23198 2428 23204 2440
rect 23159 2400 23204 2428
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 24302 2360 24308 2372
rect 22066 2332 24308 2360
rect 19116 2320 19122 2332
rect 24302 2320 24308 2332
rect 24360 2320 24366 2372
rect 24412 2360 24440 2391
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24912 2400 25145 2428
rect 24912 2388 24918 2400
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2428 25927 2431
rect 26878 2428 26884 2440
rect 25915 2400 26884 2428
rect 25915 2397 25927 2400
rect 25869 2391 25927 2397
rect 26878 2388 26884 2400
rect 26936 2388 26942 2440
rect 26988 2437 27016 2536
rect 30834 2524 30840 2536
rect 30892 2524 30898 2576
rect 32950 2524 32956 2576
rect 33008 2564 33014 2576
rect 33008 2536 35020 2564
rect 33008 2524 33014 2536
rect 30282 2496 30288 2508
rect 28092 2468 30288 2496
rect 28092 2437 28120 2468
rect 30282 2456 30288 2468
rect 30340 2456 30346 2508
rect 31478 2456 31484 2508
rect 31536 2496 31542 2508
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 31536 2468 32413 2496
rect 31536 2456 31542 2468
rect 32401 2465 32413 2468
rect 32447 2465 32459 2499
rect 32401 2459 32459 2465
rect 33318 2456 33324 2508
rect 33376 2496 33382 2508
rect 34992 2505 35020 2536
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33376 2468 34713 2496
rect 33376 2456 33382 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 34977 2499 35035 2505
rect 34977 2465 34989 2499
rect 35023 2465 35035 2499
rect 35084 2496 35112 2604
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 40405 2635 40463 2641
rect 40405 2632 40417 2635
rect 35676 2604 40417 2632
rect 35676 2592 35682 2604
rect 40405 2601 40417 2604
rect 40451 2601 40463 2635
rect 40405 2595 40463 2601
rect 45922 2592 45928 2644
rect 45980 2632 45986 2644
rect 46017 2635 46075 2641
rect 46017 2632 46029 2635
rect 45980 2604 46029 2632
rect 45980 2592 45986 2604
rect 46017 2601 46029 2604
rect 46063 2601 46075 2635
rect 46017 2595 46075 2601
rect 36998 2524 37004 2576
rect 37056 2564 37062 2576
rect 43073 2567 43131 2573
rect 43073 2564 43085 2567
rect 37056 2536 43085 2564
rect 37056 2524 37062 2536
rect 43073 2533 43085 2536
rect 43119 2533 43131 2567
rect 43073 2527 43131 2533
rect 49050 2524 49056 2576
rect 49108 2564 49114 2576
rect 49108 2536 52684 2564
rect 49108 2524 49114 2536
rect 52656 2508 52684 2536
rect 41233 2499 41291 2505
rect 41233 2496 41245 2499
rect 35084 2468 41245 2496
rect 34977 2459 35035 2465
rect 41233 2465 41245 2468
rect 41279 2465 41291 2499
rect 41233 2459 41291 2465
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 46753 2499 46811 2505
rect 46753 2496 46765 2499
rect 41380 2468 46765 2496
rect 41380 2456 41386 2468
rect 46753 2465 46765 2468
rect 46799 2465 46811 2499
rect 51258 2496 51264 2508
rect 51219 2468 51264 2496
rect 46753 2459 46811 2465
rect 51258 2456 51264 2468
rect 51316 2456 51322 2508
rect 52638 2456 52644 2508
rect 52696 2496 52702 2508
rect 52696 2468 57928 2496
rect 52696 2456 52702 2468
rect 26973 2431 27031 2437
rect 26973 2397 26985 2431
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28077 2431 28135 2437
rect 28077 2397 28089 2431
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28258 2388 28264 2440
rect 28316 2388 28322 2440
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 28960 2400 29009 2428
rect 28960 2388 28966 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 29546 2428 29552 2440
rect 29507 2400 29552 2428
rect 28997 2391 29055 2397
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 30432 2400 30481 2428
rect 30432 2388 30438 2400
rect 30469 2397 30481 2400
rect 30515 2397 30527 2431
rect 30926 2428 30932 2440
rect 30887 2400 30932 2428
rect 30469 2391 30527 2397
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 31846 2388 31852 2440
rect 31904 2428 31910 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31904 2400 32137 2428
rect 31904 2388 31910 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 33873 2431 33931 2437
rect 33873 2397 33885 2431
rect 33919 2428 33931 2431
rect 34422 2428 34428 2440
rect 33919 2400 34428 2428
rect 33919 2397 33931 2400
rect 33873 2391 33931 2397
rect 34422 2388 34428 2400
rect 34480 2388 34486 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35866 2400 36001 2428
rect 28276 2360 28304 2388
rect 24412 2332 28304 2360
rect 34698 2320 34704 2372
rect 34756 2360 34762 2372
rect 35866 2360 35894 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36262 2388 36268 2440
rect 36320 2428 36326 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36320 2400 37289 2428
rect 36320 2388 36326 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37550 2428 37556 2440
rect 37511 2400 37556 2428
rect 37277 2391 37335 2397
rect 37550 2388 37556 2400
rect 37608 2388 37614 2440
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 37660 2400 43913 2428
rect 34756 2332 35894 2360
rect 34756 2320 34762 2332
rect 37090 2320 37096 2372
rect 37148 2360 37154 2372
rect 37660 2360 37688 2400
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 45370 2388 45376 2440
rect 45428 2428 45434 2440
rect 45465 2431 45523 2437
rect 45465 2428 45477 2431
rect 45428 2400 45477 2428
rect 45428 2388 45434 2400
rect 45465 2397 45477 2400
rect 45511 2397 45523 2431
rect 45646 2428 45652 2440
rect 45607 2400 45652 2428
rect 45465 2391 45523 2397
rect 45646 2388 45652 2400
rect 45704 2388 45710 2440
rect 45830 2428 45836 2440
rect 45791 2400 45836 2428
rect 45830 2388 45836 2400
rect 45888 2388 45894 2440
rect 47946 2388 47952 2440
rect 48004 2428 48010 2440
rect 48777 2431 48835 2437
rect 48777 2428 48789 2431
rect 48004 2400 48789 2428
rect 48004 2388 48010 2400
rect 48777 2397 48789 2400
rect 48823 2397 48835 2431
rect 48777 2391 48835 2397
rect 49418 2388 49424 2440
rect 49476 2428 49482 2440
rect 50157 2431 50215 2437
rect 50157 2428 50169 2431
rect 49476 2400 50169 2428
rect 49476 2388 49482 2400
rect 50157 2397 50169 2400
rect 50203 2397 50215 2431
rect 50157 2391 50215 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 51077 2431 51135 2437
rect 51077 2428 51089 2431
rect 50948 2400 51089 2428
rect 50948 2388 50954 2400
rect 51077 2397 51089 2400
rect 51123 2397 51135 2431
rect 51077 2391 51135 2397
rect 52362 2388 52368 2440
rect 52420 2428 52426 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52420 2400 52745 2428
rect 52420 2388 52426 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53834 2388 53840 2440
rect 53892 2428 53898 2440
rect 53929 2431 53987 2437
rect 53929 2428 53941 2431
rect 53892 2400 53941 2428
rect 53892 2388 53898 2400
rect 53929 2397 53941 2400
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 55272 2400 55321 2428
rect 55272 2388 55278 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 56686 2388 56692 2440
rect 56744 2428 56750 2440
rect 57900 2437 57928 2468
rect 56781 2431 56839 2437
rect 56781 2428 56793 2431
rect 56744 2400 56793 2428
rect 56744 2388 56750 2400
rect 56781 2397 56793 2400
rect 56827 2397 56839 2431
rect 56781 2391 56839 2397
rect 57885 2431 57943 2437
rect 57885 2397 57897 2431
rect 57931 2397 57943 2431
rect 57885 2391 57943 2397
rect 37148 2332 37688 2360
rect 37148 2320 37154 2332
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 38657 2363 38715 2369
rect 38657 2360 38669 2363
rect 37792 2332 38669 2360
rect 37792 2320 37798 2332
rect 38657 2329 38669 2332
rect 38703 2329 38715 2363
rect 38657 2323 38715 2329
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39264 2332 40325 2360
rect 39264 2320 39270 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41049 2363 41107 2369
rect 41049 2360 41061 2363
rect 40644 2332 41061 2360
rect 40644 2320 40650 2332
rect 41049 2329 41061 2332
rect 41095 2329 41107 2363
rect 41049 2323 41107 2329
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 42116 2332 42901 2360
rect 42116 2320 42122 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42889 2323 42947 2329
rect 43530 2320 43536 2372
rect 43588 2360 43594 2372
rect 43717 2363 43775 2369
rect 43717 2360 43729 2363
rect 43588 2332 43729 2360
rect 43588 2320 43594 2332
rect 43717 2329 43729 2332
rect 43763 2329 43775 2363
rect 45738 2360 45744 2372
rect 45699 2332 45744 2360
rect 43717 2323 43775 2329
rect 45738 2320 45744 2332
rect 45796 2320 45802 2372
rect 46569 2363 46627 2369
rect 46569 2329 46581 2363
rect 46615 2329 46627 2363
rect 46569 2323 46627 2329
rect 16025 2295 16083 2301
rect 16025 2292 16037 2295
rect 15436 2264 16037 2292
rect 15436 2252 15442 2264
rect 16025 2261 16037 2264
rect 16071 2261 16083 2295
rect 16025 2255 16083 2261
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2261 18659 2295
rect 18601 2255 18659 2261
rect 19150 2252 19156 2304
rect 19208 2292 19214 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19208 2264 19441 2292
rect 19208 2252 19214 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20036 2264 20177 2292
rect 20036 2252 20042 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20530 2252 20536 2304
rect 20588 2292 20594 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20588 2264 20913 2292
rect 20588 2252 20594 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 24728 2264 25329 2292
rect 24728 2252 24734 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 26510 2252 26516 2304
rect 26568 2292 26574 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26568 2264 27169 2292
rect 26568 2252 26574 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 27982 2252 27988 2304
rect 28040 2292 28046 2304
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 28040 2264 28273 2292
rect 28040 2252 28046 2264
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 29454 2252 29460 2304
rect 29512 2292 29518 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 29512 2264 29745 2292
rect 29512 2252 29518 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 30834 2252 30840 2304
rect 30892 2292 30898 2304
rect 31113 2295 31171 2301
rect 31113 2292 31125 2295
rect 30892 2264 31125 2292
rect 30892 2252 30898 2264
rect 31113 2261 31125 2264
rect 31159 2261 31171 2295
rect 31113 2255 31171 2261
rect 33778 2252 33784 2304
rect 33836 2292 33842 2304
rect 34057 2295 34115 2301
rect 34057 2292 34069 2295
rect 33836 2264 34069 2292
rect 33836 2252 33842 2264
rect 34057 2261 34069 2264
rect 34103 2261 34115 2295
rect 34057 2255 34115 2261
rect 35250 2252 35256 2304
rect 35308 2292 35314 2304
rect 36173 2295 36231 2301
rect 36173 2292 36185 2295
rect 35308 2264 36185 2292
rect 35308 2252 35314 2264
rect 36173 2261 36185 2264
rect 36219 2261 36231 2295
rect 36173 2255 36231 2261
rect 36538 2252 36544 2304
rect 36596 2292 36602 2304
rect 37826 2292 37832 2304
rect 36596 2264 37832 2292
rect 36596 2252 36602 2264
rect 37826 2252 37832 2264
rect 37884 2252 37890 2304
rect 38746 2292 38752 2304
rect 38707 2264 38752 2292
rect 38746 2252 38752 2264
rect 38804 2252 38810 2304
rect 45002 2252 45008 2304
rect 45060 2292 45066 2304
rect 46584 2292 46612 2323
rect 46750 2320 46756 2372
rect 46808 2360 46814 2372
rect 48041 2363 48099 2369
rect 48041 2360 48053 2363
rect 46808 2332 48053 2360
rect 46808 2320 46814 2332
rect 48041 2329 48053 2332
rect 48087 2329 48099 2363
rect 48041 2323 48099 2329
rect 48222 2320 48228 2372
rect 48280 2360 48286 2372
rect 50433 2363 50491 2369
rect 50433 2360 50445 2363
rect 48280 2332 50445 2360
rect 48280 2320 48286 2332
rect 50433 2329 50445 2332
rect 50479 2329 50491 2363
rect 53006 2360 53012 2372
rect 52967 2332 53012 2360
rect 50433 2323 50491 2329
rect 53006 2320 53012 2332
rect 53064 2320 53070 2372
rect 54202 2360 54208 2372
rect 54163 2332 54208 2360
rect 54202 2320 54208 2332
rect 54260 2320 54266 2372
rect 55582 2360 55588 2372
rect 55543 2332 55588 2360
rect 55582 2320 55588 2332
rect 55640 2320 55646 2372
rect 57054 2360 57060 2372
rect 57015 2332 57060 2360
rect 57054 2320 57060 2332
rect 57112 2320 57118 2372
rect 48130 2292 48136 2304
rect 45060 2264 46612 2292
rect 48091 2264 48136 2292
rect 45060 2252 45066 2264
rect 48130 2252 48136 2264
rect 48188 2252 48194 2304
rect 48866 2292 48872 2304
rect 48827 2264 48872 2292
rect 48866 2252 48872 2264
rect 48924 2252 48930 2304
rect 57238 2252 57244 2304
rect 57296 2292 57302 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 57296 2264 58081 2292
rect 57296 2252 57302 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 6362 2048 6368 2100
rect 6420 2088 6426 2100
rect 23198 2088 23204 2100
rect 6420 2060 23204 2088
rect 6420 2048 6426 2060
rect 23198 2048 23204 2060
rect 23256 2048 23262 2100
rect 26878 2048 26884 2100
rect 26936 2088 26942 2100
rect 32030 2088 32036 2100
rect 26936 2060 32036 2088
rect 26936 2048 26942 2060
rect 32030 2048 32036 2060
rect 32088 2048 32094 2100
rect 37182 2048 37188 2100
rect 37240 2088 37246 2100
rect 41322 2088 41328 2100
rect 37240 2060 41328 2088
rect 37240 2048 37246 2060
rect 41322 2048 41328 2060
rect 41380 2048 41386 2100
rect 12986 1980 12992 2032
rect 13044 2020 13050 2032
rect 22002 2020 22008 2032
rect 13044 1992 22008 2020
rect 13044 1980 13050 1992
rect 22002 1980 22008 1992
rect 22060 1980 22066 2032
rect 31662 1980 31668 2032
rect 31720 2020 31726 2032
rect 37550 2020 37556 2032
rect 31720 1992 37556 2020
rect 31720 1980 31726 1992
rect 37550 1980 37556 1992
rect 37608 1980 37614 2032
rect 37826 1980 37832 2032
rect 37884 2020 37890 2032
rect 48130 2020 48136 2032
rect 37884 1992 48136 2020
rect 37884 1980 37890 1992
rect 48130 1980 48136 1992
rect 48188 1980 48194 2032
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 57054 1952 57060 1964
rect 16356 1924 57060 1952
rect 16356 1912 16362 1924
rect 57054 1912 57060 1924
rect 57112 1912 57118 1964
rect 20438 1844 20444 1896
rect 20496 1884 20502 1896
rect 45738 1884 45744 1896
rect 20496 1856 45744 1884
rect 20496 1844 20502 1856
rect 45738 1844 45744 1856
rect 45796 1844 45802 1896
rect 16390 1776 16396 1828
rect 16448 1816 16454 1828
rect 55582 1816 55588 1828
rect 16448 1788 55588 1816
rect 16448 1776 16454 1788
rect 55582 1776 55588 1788
rect 55640 1776 55646 1828
rect 12710 1708 12716 1760
rect 12768 1748 12774 1760
rect 54202 1748 54208 1760
rect 12768 1720 54208 1748
rect 12768 1708 12774 1720
rect 54202 1708 54208 1720
rect 54260 1708 54266 1760
rect 10226 1640 10232 1692
rect 10284 1680 10290 1692
rect 48222 1680 48228 1692
rect 10284 1652 48228 1680
rect 10284 1640 10290 1652
rect 48222 1640 48228 1652
rect 48280 1640 48286 1692
rect 10686 1572 10692 1624
rect 10744 1612 10750 1624
rect 53006 1612 53012 1624
rect 10744 1584 53012 1612
rect 10744 1572 10750 1584
rect 53006 1572 53012 1584
rect 53064 1572 53070 1624
rect 37642 1504 37648 1556
rect 37700 1544 37706 1556
rect 48866 1544 48872 1556
rect 37700 1516 48872 1544
rect 37700 1504 37706 1516
rect 48866 1504 48872 1516
rect 48924 1504 48930 1556
rect 7098 1436 7104 1488
rect 7156 1476 7162 1488
rect 22738 1476 22744 1488
rect 7156 1448 22744 1476
rect 7156 1436 7162 1448
rect 22738 1436 22744 1448
rect 22796 1436 22802 1488
rect 33502 1436 33508 1488
rect 33560 1476 33566 1488
rect 38746 1476 38752 1488
rect 33560 1448 38752 1476
rect 33560 1436 33566 1448
rect 38746 1436 38752 1448
rect 38804 1436 38810 1488
rect 3326 1028 3332 1080
rect 3384 1068 3390 1080
rect 8570 1068 8576 1080
rect 3384 1040 8576 1068
rect 3384 1028 3390 1040
rect 8570 1028 8576 1040
rect 8628 1028 8634 1080
<< via1 >>
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2780 39584 2832 39636
rect 3056 39627 3108 39636
rect 3056 39593 3065 39627
rect 3065 39593 3099 39627
rect 3099 39593 3108 39627
rect 3056 39584 3108 39593
rect 3700 39584 3752 39636
rect 26240 39584 26292 39636
rect 41420 39627 41472 39636
rect 41420 39593 41429 39627
rect 41429 39593 41463 39627
rect 41463 39593 41472 39627
rect 41420 39584 41472 39593
rect 48688 39584 48740 39636
rect 56140 39584 56192 39636
rect 18696 39448 18748 39500
rect 1768 39380 1820 39432
rect 2320 39380 2372 39432
rect 2872 39423 2924 39432
rect 2872 39389 2881 39423
rect 2881 39389 2915 39423
rect 2915 39389 2924 39423
rect 2872 39380 2924 39389
rect 4068 39380 4120 39432
rect 32128 39380 32180 39432
rect 33692 39380 33744 39432
rect 54760 39380 54812 39432
rect 1584 39287 1636 39296
rect 1584 39253 1593 39287
rect 1593 39253 1627 39287
rect 1627 39253 1636 39287
rect 1584 39244 1636 39253
rect 43444 39244 43496 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 32128 39083 32180 39092
rect 32128 39049 32137 39083
rect 32137 39049 32171 39083
rect 32171 39049 32180 39083
rect 32128 39040 32180 39049
rect 13268 38904 13320 38956
rect 32496 38904 32548 38956
rect 1584 38743 1636 38752
rect 1584 38709 1593 38743
rect 1593 38709 1627 38743
rect 1627 38709 1636 38743
rect 1584 38700 1636 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2964 38496 3016 38548
rect 14464 38292 14516 38344
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 1676 37816 1728 37868
rect 1584 37655 1636 37664
rect 1584 37621 1593 37655
rect 1593 37621 1627 37655
rect 1627 37621 1636 37655
rect 1584 37612 1636 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 12072 36728 12124 36780
rect 1584 36635 1636 36644
rect 1584 36601 1593 36635
rect 1593 36601 1627 36635
rect 1627 36601 1636 36635
rect 1584 36592 1636 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2044 36116 2096 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1860 35003 1912 35012
rect 1860 34969 1869 35003
rect 1869 34969 1903 35003
rect 1903 34969 1912 35003
rect 1860 34960 1912 34969
rect 1952 34935 2004 34944
rect 1952 34901 1961 34935
rect 1961 34901 1995 34935
rect 1995 34901 2004 34935
rect 1952 34892 2004 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 1584 34731 1636 34740
rect 1584 34697 1593 34731
rect 1593 34697 1627 34731
rect 1627 34697 1636 34731
rect 1584 34688 1636 34697
rect 6552 34688 6604 34740
rect 2320 34595 2372 34604
rect 2320 34561 2329 34595
rect 2329 34561 2363 34595
rect 2363 34561 2372 34595
rect 2320 34552 2372 34561
rect 6184 34484 6236 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9496 33940 9548 33992
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 2780 33464 2832 33516
rect 2228 33396 2280 33448
rect 6644 33260 6696 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17040 32852 17092 32904
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 21916 32172 21968 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4988 31968 5040 32020
rect 15476 31900 15528 31952
rect 2320 31807 2372 31816
rect 2320 31773 2329 31807
rect 2329 31773 2363 31807
rect 2363 31773 2372 31807
rect 2320 31764 2372 31773
rect 1584 31671 1636 31680
rect 1584 31637 1593 31671
rect 1593 31637 1627 31671
rect 1627 31637 1636 31671
rect 1584 31628 1636 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 1768 31331 1820 31340
rect 1768 31297 1777 31331
rect 1777 31297 1811 31331
rect 1811 31297 1820 31331
rect 1768 31288 1820 31297
rect 2504 31263 2556 31272
rect 2504 31229 2513 31263
rect 2513 31229 2547 31263
rect 2547 31229 2556 31263
rect 2504 31220 2556 31229
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 12900 30744 12952 30796
rect 2412 30719 2464 30728
rect 2412 30685 2421 30719
rect 2421 30685 2455 30719
rect 2455 30685 2464 30719
rect 2412 30676 2464 30685
rect 3056 30719 3108 30728
rect 3056 30685 3065 30719
rect 3065 30685 3099 30719
rect 3099 30685 3108 30719
rect 3056 30676 3108 30685
rect 4896 30719 4948 30728
rect 4896 30685 4905 30719
rect 4905 30685 4939 30719
rect 4939 30685 4948 30719
rect 4896 30676 4948 30685
rect 1584 30583 1636 30592
rect 1584 30549 1593 30583
rect 1593 30549 1627 30583
rect 1627 30549 1636 30583
rect 1584 30540 1636 30549
rect 2320 30540 2372 30592
rect 2688 30540 2740 30592
rect 4712 30583 4764 30592
rect 4712 30549 4721 30583
rect 4721 30549 4755 30583
rect 4755 30549 4764 30583
rect 4712 30540 4764 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4712 30311 4764 30320
rect 1400 30200 1452 30252
rect 1860 30132 1912 30184
rect 2320 30243 2372 30252
rect 2320 30209 2354 30243
rect 2354 30209 2372 30243
rect 2320 30200 2372 30209
rect 4712 30277 4746 30311
rect 4746 30277 4764 30311
rect 4712 30268 4764 30277
rect 3056 29996 3108 30048
rect 3424 30039 3476 30048
rect 3424 30005 3433 30039
rect 3433 30005 3467 30039
rect 3467 30005 3476 30039
rect 3424 29996 3476 30005
rect 5080 29996 5132 30048
rect 5816 30039 5868 30048
rect 5816 30005 5825 30039
rect 5825 30005 5859 30039
rect 5859 30005 5868 30039
rect 5816 29996 5868 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2412 29792 2464 29844
rect 4896 29792 4948 29844
rect 5080 29792 5132 29844
rect 2596 29724 2648 29776
rect 2688 29656 2740 29708
rect 4988 29699 5040 29708
rect 4988 29665 4997 29699
rect 4997 29665 5031 29699
rect 5031 29665 5040 29699
rect 4988 29656 5040 29665
rect 1676 29631 1728 29640
rect 1676 29597 1685 29631
rect 1685 29597 1719 29631
rect 1719 29597 1728 29631
rect 1676 29588 1728 29597
rect 5816 29588 5868 29640
rect 6736 29588 6788 29640
rect 3424 29520 3476 29572
rect 6368 29563 6420 29572
rect 6368 29529 6377 29563
rect 6377 29529 6411 29563
rect 6411 29529 6420 29563
rect 6368 29520 6420 29529
rect 3332 29452 3384 29504
rect 7104 29452 7156 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 1676 29248 1728 29300
rect 2136 29248 2188 29300
rect 6368 29248 6420 29300
rect 12900 29291 12952 29300
rect 12900 29257 12909 29291
rect 12909 29257 12943 29291
rect 12943 29257 12952 29291
rect 12900 29248 12952 29257
rect 15476 29291 15528 29300
rect 15476 29257 15485 29291
rect 15485 29257 15519 29291
rect 15519 29257 15528 29291
rect 15476 29248 15528 29257
rect 2688 29112 2740 29164
rect 2872 29112 2924 29164
rect 5816 29155 5868 29164
rect 5816 29121 5825 29155
rect 5825 29121 5859 29155
rect 5859 29121 5868 29155
rect 5816 29112 5868 29121
rect 12348 29180 12400 29232
rect 12164 29112 12216 29164
rect 14740 29112 14792 29164
rect 1860 29044 1912 29096
rect 2136 29044 2188 29096
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 2780 28976 2832 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2872 28704 2924 28756
rect 5816 28704 5868 28756
rect 12164 28747 12216 28756
rect 12164 28713 12173 28747
rect 12173 28713 12207 28747
rect 12207 28713 12216 28747
rect 12164 28704 12216 28713
rect 14740 28747 14792 28756
rect 14740 28713 14749 28747
rect 14749 28713 14783 28747
rect 14783 28713 14792 28747
rect 14740 28704 14792 28713
rect 2596 28568 2648 28620
rect 6644 28611 6696 28620
rect 6644 28577 6653 28611
rect 6653 28577 6687 28611
rect 6687 28577 6696 28611
rect 6644 28568 6696 28577
rect 6828 28611 6880 28620
rect 6828 28577 6837 28611
rect 6837 28577 6871 28611
rect 6871 28577 6880 28611
rect 6828 28568 6880 28577
rect 6368 28500 6420 28552
rect 12624 28543 12676 28552
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 3056 28432 3108 28484
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 12624 28500 12676 28509
rect 1768 28364 1820 28416
rect 3884 28364 3936 28416
rect 6736 28364 6788 28416
rect 7288 28364 7340 28416
rect 12900 28432 12952 28484
rect 13728 28364 13780 28416
rect 17132 28500 17184 28552
rect 17316 28543 17368 28552
rect 17316 28509 17325 28543
rect 17325 28509 17359 28543
rect 17359 28509 17368 28543
rect 17316 28500 17368 28509
rect 15476 28432 15528 28484
rect 18052 28432 18104 28484
rect 16580 28364 16632 28416
rect 18696 28407 18748 28416
rect 18696 28373 18705 28407
rect 18705 28373 18739 28407
rect 18739 28373 18748 28407
rect 18696 28364 18748 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2688 28160 2740 28212
rect 17040 28203 17092 28212
rect 2780 28135 2832 28144
rect 2780 28101 2814 28135
rect 2814 28101 2832 28135
rect 2780 28092 2832 28101
rect 17040 28169 17049 28203
rect 17049 28169 17083 28203
rect 17083 28169 17092 28203
rect 17040 28160 17092 28169
rect 18052 28203 18104 28212
rect 18052 28169 18061 28203
rect 18061 28169 18095 28203
rect 18095 28169 18104 28203
rect 18052 28160 18104 28169
rect 18696 28092 18748 28144
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 17132 28024 17184 28033
rect 18236 28067 18288 28076
rect 18236 28033 18245 28067
rect 18245 28033 18279 28067
rect 18279 28033 18288 28067
rect 18236 28024 18288 28033
rect 2136 27956 2188 28008
rect 18696 27956 18748 28008
rect 3884 27931 3936 27940
rect 3884 27897 3893 27931
rect 3893 27897 3927 27931
rect 3927 27897 3936 27931
rect 3884 27888 3936 27897
rect 6736 27888 6788 27940
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 16672 27863 16724 27872
rect 16672 27829 16681 27863
rect 16681 27829 16715 27863
rect 16715 27829 16724 27863
rect 16672 27820 16724 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 17040 27616 17092 27668
rect 2320 27548 2372 27600
rect 5816 27548 5868 27600
rect 2320 27412 2372 27464
rect 3976 27455 4028 27464
rect 3976 27421 3985 27455
rect 3985 27421 4019 27455
rect 4019 27421 4028 27455
rect 3976 27412 4028 27421
rect 5356 27455 5408 27464
rect 5356 27421 5365 27455
rect 5365 27421 5399 27455
rect 5399 27421 5408 27455
rect 5356 27412 5408 27421
rect 5724 27412 5776 27464
rect 9588 27412 9640 27464
rect 12348 27480 12400 27532
rect 15292 27523 15344 27532
rect 15292 27489 15301 27523
rect 15301 27489 15335 27523
rect 15335 27489 15344 27523
rect 15292 27480 15344 27489
rect 1860 27387 1912 27396
rect 1860 27353 1869 27387
rect 1869 27353 1903 27387
rect 1903 27353 1912 27387
rect 1860 27344 1912 27353
rect 2688 27319 2740 27328
rect 2688 27285 2697 27319
rect 2697 27285 2731 27319
rect 2731 27285 2740 27319
rect 2688 27276 2740 27285
rect 2780 27276 2832 27328
rect 6184 27344 6236 27396
rect 6644 27276 6696 27328
rect 10508 27344 10560 27396
rect 10876 27276 10928 27328
rect 16672 27412 16724 27464
rect 25504 27344 25556 27396
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1400 27072 1452 27124
rect 2688 27004 2740 27056
rect 5356 27072 5408 27124
rect 6552 27072 6604 27124
rect 9496 27072 9548 27124
rect 10508 27115 10560 27124
rect 10508 27081 10517 27115
rect 10517 27081 10551 27115
rect 10551 27081 10560 27115
rect 10508 27072 10560 27081
rect 10876 27115 10928 27124
rect 10876 27081 10885 27115
rect 10885 27081 10919 27115
rect 10919 27081 10928 27115
rect 10876 27072 10928 27081
rect 14464 27072 14516 27124
rect 3976 26979 4028 26988
rect 3976 26945 3985 26979
rect 3985 26945 4019 26979
rect 4019 26945 4028 26979
rect 3976 26936 4028 26945
rect 6644 26936 6696 26988
rect 9036 26936 9088 26988
rect 1400 26868 1452 26920
rect 6828 26868 6880 26920
rect 3332 26843 3384 26852
rect 3332 26809 3341 26843
rect 3341 26809 3375 26843
rect 3375 26809 3384 26843
rect 3332 26800 3384 26809
rect 5908 26800 5960 26852
rect 2136 26732 2188 26784
rect 4988 26732 5040 26784
rect 6184 26732 6236 26784
rect 13176 27004 13228 27056
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 12348 26936 12400 26988
rect 14740 26936 14792 26988
rect 15292 26936 15344 26988
rect 17316 26936 17368 26988
rect 18144 26979 18196 26988
rect 18144 26945 18178 26979
rect 18178 26945 18196 26979
rect 18144 26936 18196 26945
rect 18604 26732 18656 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2320 26571 2372 26580
rect 2320 26537 2329 26571
rect 2329 26537 2363 26571
rect 2363 26537 2372 26571
rect 2320 26528 2372 26537
rect 2596 26460 2648 26512
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 2780 26392 2832 26401
rect 5724 26528 5776 26580
rect 6184 26528 6236 26580
rect 9036 26528 9088 26580
rect 12624 26528 12676 26580
rect 14740 26571 14792 26580
rect 14740 26537 14749 26571
rect 14749 26537 14783 26571
rect 14783 26537 14792 26571
rect 14740 26528 14792 26537
rect 6000 26460 6052 26512
rect 16764 26528 16816 26580
rect 18144 26528 18196 26580
rect 4528 26367 4580 26376
rect 3332 26256 3384 26308
rect 4528 26333 4537 26367
rect 4537 26333 4571 26367
rect 4571 26333 4580 26367
rect 4528 26324 4580 26333
rect 14004 26392 14056 26444
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 9496 26367 9548 26376
rect 9496 26333 9505 26367
rect 9505 26333 9539 26367
rect 9539 26333 9548 26367
rect 9496 26324 9548 26333
rect 10140 26324 10192 26376
rect 10968 26324 11020 26376
rect 14464 26367 14516 26376
rect 12348 26299 12400 26308
rect 12348 26265 12357 26299
rect 12357 26265 12391 26299
rect 12391 26265 12400 26299
rect 12348 26256 12400 26265
rect 14464 26333 14473 26367
rect 14473 26333 14507 26367
rect 14507 26333 14516 26367
rect 14464 26324 14516 26333
rect 14556 26367 14608 26376
rect 14556 26333 14570 26367
rect 14570 26333 14604 26367
rect 14604 26333 14608 26367
rect 14556 26324 14608 26333
rect 15292 26392 15344 26444
rect 18420 26367 18472 26376
rect 18420 26333 18429 26367
rect 18429 26333 18463 26367
rect 18463 26333 18472 26367
rect 18420 26324 18472 26333
rect 18604 26367 18656 26376
rect 18604 26333 18613 26367
rect 18613 26333 18647 26367
rect 18647 26333 18656 26367
rect 18604 26324 18656 26333
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 14372 26299 14424 26308
rect 14372 26265 14381 26299
rect 14381 26265 14415 26299
rect 14415 26265 14424 26299
rect 14372 26256 14424 26265
rect 14924 26256 14976 26308
rect 16212 26256 16264 26308
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 6368 26231 6420 26240
rect 6368 26197 6377 26231
rect 6377 26197 6411 26231
rect 6411 26197 6420 26231
rect 6368 26188 6420 26197
rect 14096 26188 14148 26240
rect 15200 26188 15252 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 2596 25984 2648 26036
rect 4528 26027 4580 26036
rect 4528 25993 4537 26027
rect 4537 25993 4571 26027
rect 4571 25993 4580 26027
rect 4528 25984 4580 25993
rect 4988 26027 5040 26036
rect 4988 25993 4997 26027
rect 4997 25993 5031 26027
rect 5031 25993 5040 26027
rect 4988 25984 5040 25993
rect 16212 25984 16264 26036
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 4620 25848 4672 25900
rect 5724 25916 5776 25968
rect 6368 25916 6420 25968
rect 14372 25916 14424 25968
rect 12440 25848 12492 25900
rect 14740 25848 14792 25900
rect 15200 25848 15252 25900
rect 16764 25916 16816 25968
rect 15936 25891 15988 25900
rect 15936 25857 15950 25891
rect 15950 25857 15984 25891
rect 15984 25857 15988 25891
rect 15936 25848 15988 25857
rect 16396 25780 16448 25832
rect 5448 25712 5500 25764
rect 2136 25687 2188 25696
rect 2136 25653 2145 25687
rect 2145 25653 2179 25687
rect 2179 25653 2188 25687
rect 2136 25644 2188 25653
rect 2964 25644 3016 25696
rect 14464 25644 14516 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2136 25440 2188 25492
rect 27068 25440 27120 25492
rect 14740 25415 14792 25424
rect 14740 25381 14749 25415
rect 14749 25381 14783 25415
rect 14783 25381 14792 25415
rect 14740 25372 14792 25381
rect 2320 25236 2372 25288
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 8852 25236 8904 25288
rect 9588 25236 9640 25288
rect 12440 25236 12492 25288
rect 14096 25279 14148 25288
rect 14096 25245 14105 25279
rect 14105 25245 14139 25279
rect 14139 25245 14148 25279
rect 14096 25236 14148 25245
rect 14464 25279 14516 25288
rect 4620 25168 4672 25220
rect 10232 25168 10284 25220
rect 11060 25211 11112 25220
rect 11060 25177 11094 25211
rect 11094 25177 11112 25211
rect 11060 25168 11112 25177
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 2412 25100 2464 25152
rect 6276 25100 6328 25152
rect 6828 25100 6880 25152
rect 9864 25100 9916 25152
rect 10048 25100 10100 25152
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 14556 25279 14608 25288
rect 14556 25245 14570 25279
rect 14570 25245 14604 25279
rect 14604 25245 14608 25279
rect 14556 25236 14608 25245
rect 14372 25211 14424 25220
rect 14372 25177 14381 25211
rect 14381 25177 14415 25211
rect 14415 25177 14424 25211
rect 14372 25168 14424 25177
rect 15016 25143 15068 25152
rect 15016 25109 15025 25143
rect 15025 25109 15059 25143
rect 15059 25109 15068 25143
rect 15016 25100 15068 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 5448 24896 5500 24948
rect 10232 24896 10284 24948
rect 1676 24828 1728 24880
rect 10048 24871 10100 24880
rect 10048 24837 10057 24871
rect 10057 24837 10091 24871
rect 10091 24837 10100 24871
rect 10048 24828 10100 24837
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 1400 24692 1452 24744
rect 1492 24692 1544 24744
rect 1676 24692 1728 24744
rect 2228 24760 2280 24812
rect 2412 24803 2464 24812
rect 2412 24769 2446 24803
rect 2446 24769 2464 24803
rect 2412 24760 2464 24769
rect 5172 24692 5224 24744
rect 3516 24667 3568 24676
rect 3516 24633 3525 24667
rect 3525 24633 3559 24667
rect 3559 24633 3568 24667
rect 3516 24624 3568 24633
rect 5816 24624 5868 24676
rect 1400 24599 1452 24608
rect 1400 24565 1409 24599
rect 1409 24565 1443 24599
rect 1443 24565 1452 24599
rect 1400 24556 1452 24565
rect 5632 24556 5684 24608
rect 6276 24760 6328 24812
rect 6184 24692 6236 24744
rect 9772 24803 9824 24812
rect 9772 24769 9782 24803
rect 9782 24769 9816 24803
rect 9816 24769 9824 24803
rect 9772 24760 9824 24769
rect 10140 24803 10192 24812
rect 10140 24769 10154 24803
rect 10154 24769 10188 24803
rect 10188 24769 10192 24803
rect 10140 24760 10192 24769
rect 13636 24760 13688 24812
rect 14556 24760 14608 24812
rect 15660 24760 15712 24812
rect 15936 24760 15988 24812
rect 18328 24760 18380 24812
rect 10600 24692 10652 24744
rect 15476 24692 15528 24744
rect 18880 24735 18932 24744
rect 18880 24701 18889 24735
rect 18889 24701 18923 24735
rect 18923 24701 18932 24735
rect 18880 24692 18932 24701
rect 10324 24624 10376 24676
rect 6368 24556 6420 24608
rect 14004 24556 14056 24608
rect 18604 24556 18656 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2504 24352 2556 24404
rect 6184 24352 6236 24404
rect 8852 24352 8904 24404
rect 11060 24352 11112 24404
rect 18328 24352 18380 24404
rect 2412 24284 2464 24336
rect 1400 24216 1452 24268
rect 10324 24284 10376 24336
rect 5172 24259 5224 24268
rect 5172 24225 5181 24259
rect 5181 24225 5215 24259
rect 5215 24225 5224 24259
rect 5172 24216 5224 24225
rect 10140 24216 10192 24268
rect 1492 24191 1544 24200
rect 1492 24157 1501 24191
rect 1501 24157 1535 24191
rect 1535 24157 1544 24191
rect 1492 24148 1544 24157
rect 3516 24148 3568 24200
rect 1676 24080 1728 24132
rect 10232 24148 10284 24200
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10508 24191 10560 24200
rect 10324 24148 10376 24157
rect 10508 24157 10515 24191
rect 10515 24157 10560 24191
rect 10508 24148 10560 24157
rect 12532 24216 12584 24268
rect 15476 24216 15528 24268
rect 18880 24216 18932 24268
rect 12716 24148 12768 24200
rect 13268 24191 13320 24200
rect 4620 24080 4672 24132
rect 10600 24123 10652 24132
rect 10600 24089 10609 24123
rect 10609 24089 10643 24123
rect 10643 24089 10652 24123
rect 10600 24080 10652 24089
rect 12164 24080 12216 24132
rect 12808 24080 12860 24132
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 13636 24148 13688 24200
rect 18696 24191 18748 24200
rect 14372 24080 14424 24132
rect 15844 24123 15896 24132
rect 15844 24089 15878 24123
rect 15878 24089 15896 24123
rect 15844 24080 15896 24089
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 2044 24012 2096 24064
rect 13360 24012 13412 24064
rect 13544 24055 13596 24064
rect 13544 24021 13553 24055
rect 13553 24021 13587 24055
rect 13587 24021 13596 24055
rect 13544 24012 13596 24021
rect 16948 24055 17000 24064
rect 16948 24021 16957 24055
rect 16957 24021 16991 24055
rect 16991 24021 17000 24055
rect 16948 24012 17000 24021
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 18604 24123 18656 24132
rect 18604 24089 18613 24123
rect 18613 24089 18647 24123
rect 18647 24089 18656 24123
rect 18604 24080 18656 24089
rect 19064 24080 19116 24132
rect 20260 24012 20312 24064
rect 20628 24055 20680 24064
rect 20628 24021 20637 24055
rect 20637 24021 20671 24055
rect 20671 24021 20680 24055
rect 20628 24012 20680 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 2320 23808 2372 23860
rect 2596 23740 2648 23792
rect 6368 23783 6420 23792
rect 6368 23749 6377 23783
rect 6377 23749 6411 23783
rect 6411 23749 6420 23783
rect 6368 23740 6420 23749
rect 6920 23740 6972 23792
rect 10140 23740 10192 23792
rect 2228 23672 2280 23724
rect 2688 23672 2740 23724
rect 5080 23672 5132 23724
rect 7196 23672 7248 23724
rect 10416 23672 10468 23724
rect 12072 23672 12124 23724
rect 13360 23808 13412 23860
rect 15844 23851 15896 23860
rect 13544 23740 13596 23792
rect 14372 23740 14424 23792
rect 14832 23740 14884 23792
rect 15844 23817 15853 23851
rect 15853 23817 15887 23851
rect 15887 23817 15896 23851
rect 15844 23808 15896 23817
rect 19064 23851 19116 23860
rect 19064 23817 19073 23851
rect 19073 23817 19107 23851
rect 19107 23817 19116 23851
rect 19064 23808 19116 23817
rect 16948 23740 17000 23792
rect 5816 23604 5868 23656
rect 8852 23647 8904 23656
rect 8852 23613 8861 23647
rect 8861 23613 8895 23647
rect 8895 23613 8904 23647
rect 8852 23604 8904 23613
rect 12440 23604 12492 23656
rect 1768 23468 1820 23520
rect 2044 23468 2096 23520
rect 3516 23511 3568 23520
rect 3516 23477 3525 23511
rect 3525 23477 3559 23511
rect 3559 23477 3568 23511
rect 3516 23468 3568 23477
rect 6368 23511 6420 23520
rect 6368 23477 6377 23511
rect 6377 23477 6411 23511
rect 6411 23477 6420 23511
rect 6368 23468 6420 23477
rect 7472 23468 7524 23520
rect 10232 23579 10284 23588
rect 10232 23545 10241 23579
rect 10241 23545 10275 23579
rect 10275 23545 10284 23579
rect 10232 23536 10284 23545
rect 9588 23468 9640 23520
rect 15200 23715 15252 23724
rect 15200 23681 15209 23715
rect 15209 23681 15243 23715
rect 15243 23681 15252 23715
rect 15200 23672 15252 23681
rect 15660 23715 15712 23724
rect 20536 23808 20588 23860
rect 20628 23740 20680 23792
rect 15660 23681 15674 23715
rect 15674 23681 15708 23715
rect 15708 23681 15712 23715
rect 15660 23672 15712 23681
rect 16488 23604 16540 23656
rect 12992 23468 13044 23520
rect 13452 23468 13504 23520
rect 15200 23468 15252 23520
rect 15752 23468 15804 23520
rect 18696 23468 18748 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2688 23307 2740 23316
rect 2688 23273 2697 23307
rect 2697 23273 2731 23307
rect 2731 23273 2740 23307
rect 2688 23264 2740 23273
rect 5816 23307 5868 23316
rect 5816 23273 5825 23307
rect 5825 23273 5859 23307
rect 5859 23273 5868 23307
rect 5816 23264 5868 23273
rect 5908 23264 5960 23316
rect 10416 23307 10468 23316
rect 10416 23273 10425 23307
rect 10425 23273 10459 23307
rect 10459 23273 10468 23307
rect 10416 23264 10468 23273
rect 14832 23307 14884 23316
rect 14832 23273 14841 23307
rect 14841 23273 14875 23307
rect 14875 23273 14884 23307
rect 14832 23264 14884 23273
rect 7656 23196 7708 23248
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 5724 23171 5776 23180
rect 5724 23137 5733 23171
rect 5733 23137 5767 23171
rect 5767 23137 5776 23171
rect 6644 23171 6696 23180
rect 5724 23128 5776 23137
rect 1676 23103 1728 23112
rect 1676 23069 1685 23103
rect 1685 23069 1719 23103
rect 1719 23069 1728 23103
rect 1676 23060 1728 23069
rect 2228 23060 2280 23112
rect 3976 23103 4028 23112
rect 3976 23069 3985 23103
rect 3985 23069 4019 23103
rect 4019 23069 4028 23103
rect 3976 23060 4028 23069
rect 3516 22992 3568 23044
rect 6368 23060 6420 23112
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 10324 23196 10376 23248
rect 13636 23196 13688 23248
rect 10048 23128 10100 23180
rect 9956 23103 10008 23112
rect 9956 23069 9963 23103
rect 9963 23069 10008 23103
rect 9956 23060 10008 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 15476 23128 15528 23180
rect 12072 23060 12124 23112
rect 14832 23060 14884 23112
rect 21640 23060 21692 23112
rect 24676 23060 24728 23112
rect 27988 23060 28040 23112
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 31208 23060 31260 23069
rect 34612 23060 34664 23112
rect 5908 22992 5960 23044
rect 7840 22992 7892 23044
rect 10324 22992 10376 23044
rect 10600 22992 10652 23044
rect 12900 22992 12952 23044
rect 16764 22992 16816 23044
rect 22100 22992 22152 23044
rect 25780 22992 25832 23044
rect 31484 23035 31536 23044
rect 31484 23001 31518 23035
rect 31518 23001 31536 23035
rect 31484 22992 31536 23001
rect 2688 22924 2740 22976
rect 7380 22924 7432 22976
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 12348 22924 12400 22976
rect 17408 22967 17460 22976
rect 17408 22933 17417 22967
rect 17417 22933 17451 22967
rect 17451 22933 17460 22967
rect 17408 22924 17460 22933
rect 21732 22924 21784 22976
rect 26792 22967 26844 22976
rect 26792 22933 26801 22967
rect 26801 22933 26835 22967
rect 26835 22933 26844 22967
rect 26792 22924 26844 22933
rect 28448 22967 28500 22976
rect 28448 22933 28457 22967
rect 28457 22933 28491 22967
rect 28491 22933 28500 22967
rect 28448 22924 28500 22933
rect 32220 22924 32272 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 2688 22763 2740 22772
rect 2688 22729 2697 22763
rect 2697 22729 2731 22763
rect 2731 22729 2740 22763
rect 2688 22720 2740 22729
rect 2780 22720 2832 22772
rect 16764 22763 16816 22772
rect 1676 22652 1728 22704
rect 13084 22652 13136 22704
rect 16764 22729 16773 22763
rect 16773 22729 16807 22763
rect 16807 22729 16816 22763
rect 16764 22720 16816 22729
rect 17408 22652 17460 22704
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 3516 22584 3568 22636
rect 3976 22627 4028 22636
rect 3976 22593 4010 22627
rect 4010 22593 4028 22627
rect 7104 22627 7156 22636
rect 3976 22584 4028 22593
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 7380 22627 7432 22636
rect 2412 22516 2464 22568
rect 2688 22516 2740 22568
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 14832 22584 14884 22636
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 18696 22720 18748 22772
rect 20352 22720 20404 22772
rect 25780 22763 25832 22772
rect 25780 22729 25789 22763
rect 25789 22729 25823 22763
rect 25823 22729 25832 22763
rect 25780 22720 25832 22729
rect 24768 22652 24820 22704
rect 26792 22720 26844 22772
rect 27988 22763 28040 22772
rect 27988 22729 27997 22763
rect 27997 22729 28031 22763
rect 28031 22729 28040 22763
rect 27988 22720 28040 22729
rect 1492 22448 1544 22500
rect 2320 22448 2372 22500
rect 7748 22516 7800 22568
rect 14280 22516 14332 22568
rect 18972 22584 19024 22636
rect 19156 22584 19208 22636
rect 19524 22627 19576 22636
rect 18604 22559 18656 22568
rect 18604 22525 18613 22559
rect 18613 22525 18647 22559
rect 18647 22525 18656 22559
rect 18604 22516 18656 22525
rect 18696 22559 18748 22568
rect 18696 22525 18705 22559
rect 18705 22525 18739 22559
rect 18739 22525 18748 22559
rect 18696 22516 18748 22525
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 5080 22423 5132 22432
rect 5080 22389 5089 22423
rect 5089 22389 5123 22423
rect 5123 22389 5132 22423
rect 5080 22380 5132 22389
rect 7012 22380 7064 22432
rect 10324 22380 10376 22432
rect 13728 22380 13780 22432
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 19524 22593 19533 22627
rect 19533 22593 19567 22627
rect 19567 22593 19576 22627
rect 19524 22584 19576 22593
rect 19800 22584 19852 22636
rect 23020 22584 23072 22636
rect 26424 22652 26476 22704
rect 28448 22652 28500 22704
rect 32220 22695 32272 22704
rect 32220 22661 32229 22695
rect 32229 22661 32263 22695
rect 32263 22661 32272 22695
rect 32220 22652 32272 22661
rect 32404 22695 32456 22704
rect 32404 22661 32429 22695
rect 32429 22661 32456 22695
rect 32404 22652 32456 22661
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 19524 22448 19576 22500
rect 21640 22516 21692 22568
rect 27896 22516 27948 22568
rect 31208 22584 31260 22636
rect 31300 22584 31352 22636
rect 32588 22584 32640 22636
rect 33140 22584 33192 22636
rect 33968 22584 34020 22636
rect 34612 22627 34664 22636
rect 34612 22593 34621 22627
rect 34621 22593 34655 22627
rect 34655 22593 34664 22627
rect 34612 22584 34664 22593
rect 34704 22584 34756 22636
rect 21732 22448 21784 22500
rect 31760 22448 31812 22500
rect 19800 22380 19852 22432
rect 23388 22380 23440 22432
rect 30196 22380 30248 22432
rect 31944 22380 31996 22432
rect 32772 22380 32824 22432
rect 34796 22380 34848 22432
rect 36268 22380 36320 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1400 22176 1452 22228
rect 2688 22108 2740 22160
rect 7104 22040 7156 22092
rect 1860 22015 1912 22024
rect 1860 21981 1869 22015
rect 1869 21981 1903 22015
rect 1903 21981 1912 22015
rect 1860 21972 1912 21981
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 5080 21972 5132 22024
rect 6644 21972 6696 22024
rect 7380 21972 7432 22024
rect 9680 22040 9732 22092
rect 10232 22040 10284 22092
rect 12992 22040 13044 22092
rect 18236 22040 18288 22092
rect 19248 22176 19300 22228
rect 20352 22219 20404 22228
rect 20352 22185 20361 22219
rect 20361 22185 20395 22219
rect 20395 22185 20404 22219
rect 20352 22176 20404 22185
rect 18604 22108 18656 22160
rect 18880 22108 18932 22160
rect 19524 22083 19576 22092
rect 19524 22049 19534 22083
rect 19534 22049 19568 22083
rect 19568 22049 19576 22083
rect 19984 22108 20036 22160
rect 19524 22040 19576 22049
rect 19800 22083 19852 22092
rect 19800 22049 19809 22083
rect 19809 22049 19843 22083
rect 19843 22049 19852 22083
rect 20812 22176 20864 22228
rect 23020 22219 23072 22228
rect 23020 22185 23029 22219
rect 23029 22185 23063 22219
rect 23063 22185 23072 22219
rect 23020 22176 23072 22185
rect 27620 22176 27672 22228
rect 28448 22176 28500 22228
rect 31484 22219 31536 22228
rect 20628 22083 20680 22092
rect 19800 22040 19852 22049
rect 20628 22049 20637 22083
rect 20637 22049 20671 22083
rect 20671 22049 20680 22083
rect 20628 22040 20680 22049
rect 23388 22108 23440 22160
rect 28816 22108 28868 22160
rect 28908 22108 28960 22160
rect 2320 21904 2372 21956
rect 7104 21904 7156 21956
rect 8208 21904 8260 21956
rect 3884 21879 3936 21888
rect 3884 21845 3893 21879
rect 3893 21845 3927 21879
rect 3927 21845 3936 21879
rect 3884 21836 3936 21845
rect 7012 21879 7064 21888
rect 7012 21845 7021 21879
rect 7021 21845 7055 21879
rect 7055 21845 7064 21879
rect 7012 21836 7064 21845
rect 7472 21836 7524 21888
rect 7748 21836 7800 21888
rect 12900 22015 12952 22024
rect 12900 21981 12909 22015
rect 12909 21981 12943 22015
rect 12943 21981 12952 22015
rect 12900 21972 12952 21981
rect 14188 21972 14240 22024
rect 13820 21904 13872 21956
rect 18696 21972 18748 22024
rect 18788 21972 18840 22024
rect 19432 21972 19484 22024
rect 20444 21972 20496 22024
rect 20812 22015 20864 22024
rect 20352 21904 20404 21956
rect 15200 21836 15252 21888
rect 15476 21879 15528 21888
rect 15476 21845 15485 21879
rect 15485 21845 15519 21879
rect 15519 21845 15528 21879
rect 15476 21836 15528 21845
rect 17868 21836 17920 21888
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 22376 21972 22428 22024
rect 22468 21972 22520 22024
rect 23112 21972 23164 22024
rect 21732 21904 21784 21956
rect 23388 21947 23440 21956
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 23020 21836 23072 21888
rect 23388 21913 23397 21947
rect 23397 21913 23431 21947
rect 23431 21913 23440 21947
rect 23388 21904 23440 21913
rect 23296 21836 23348 21888
rect 26240 21972 26292 22024
rect 31484 22185 31493 22219
rect 31493 22185 31527 22219
rect 31527 22185 31536 22219
rect 31484 22176 31536 22185
rect 34704 22219 34756 22228
rect 34704 22185 34713 22219
rect 34713 22185 34747 22219
rect 34747 22185 34756 22219
rect 34704 22176 34756 22185
rect 30196 22108 30248 22160
rect 32036 22108 32088 22160
rect 29092 21972 29144 22024
rect 30196 22015 30248 22024
rect 30196 21981 30205 22015
rect 30205 21981 30239 22015
rect 30239 21981 30248 22015
rect 30196 21972 30248 21981
rect 29184 21904 29236 21956
rect 30564 21972 30616 22024
rect 31392 21972 31444 22024
rect 31944 22015 31996 22024
rect 31944 21981 31953 22015
rect 31953 21981 31987 22015
rect 31987 21981 31996 22015
rect 31944 21972 31996 21981
rect 31484 21904 31536 21956
rect 31852 21879 31904 21888
rect 31852 21845 31861 21879
rect 31861 21845 31895 21879
rect 31895 21845 31904 21879
rect 31852 21836 31904 21845
rect 33140 22040 33192 22092
rect 32680 21972 32732 22024
rect 36268 22040 36320 22092
rect 32588 21904 32640 21956
rect 33416 22015 33468 22024
rect 33416 21981 33425 22015
rect 33425 21981 33459 22015
rect 33459 21981 33468 22015
rect 33416 21972 33468 21981
rect 33600 22015 33652 22024
rect 33600 21981 33609 22015
rect 33609 21981 33643 22015
rect 33643 21981 33652 22015
rect 33600 21972 33652 21981
rect 34796 21972 34848 22024
rect 39120 21972 39172 22024
rect 34428 21904 34480 21956
rect 37832 21904 37884 21956
rect 38292 21904 38344 21956
rect 35716 21836 35768 21888
rect 38660 21836 38712 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3976 21632 4028 21684
rect 7104 21632 7156 21684
rect 7288 21632 7340 21684
rect 7564 21632 7616 21684
rect 7748 21632 7800 21684
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 16580 21632 16632 21684
rect 18420 21632 18472 21684
rect 20444 21632 20496 21684
rect 24768 21632 24820 21684
rect 28908 21632 28960 21684
rect 15476 21564 15528 21616
rect 15568 21564 15620 21616
rect 1768 21496 1820 21548
rect 2044 21496 2096 21548
rect 2412 21539 2464 21548
rect 2412 21505 2421 21539
rect 2421 21505 2455 21539
rect 2455 21505 2464 21539
rect 2412 21496 2464 21505
rect 3056 21539 3108 21548
rect 3056 21505 3065 21539
rect 3065 21505 3099 21539
rect 3099 21505 3108 21539
rect 3056 21496 3108 21505
rect 3884 21496 3936 21548
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 7288 21496 7340 21548
rect 7748 21496 7800 21548
rect 8116 21496 8168 21548
rect 8208 21496 8260 21548
rect 14280 21539 14332 21548
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 8024 21428 8076 21480
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 2228 21335 2280 21344
rect 2228 21301 2237 21335
rect 2237 21301 2271 21335
rect 2271 21301 2280 21335
rect 2228 21292 2280 21301
rect 2872 21335 2924 21344
rect 2872 21301 2881 21335
rect 2881 21301 2915 21335
rect 2915 21301 2924 21335
rect 2872 21292 2924 21301
rect 6920 21292 6972 21344
rect 7288 21292 7340 21344
rect 7748 21292 7800 21344
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 8208 21335 8260 21344
rect 7840 21292 7892 21301
rect 8208 21301 8217 21335
rect 8217 21301 8251 21335
rect 8251 21301 8260 21335
rect 8208 21292 8260 21301
rect 14280 21505 14289 21539
rect 14289 21505 14323 21539
rect 14323 21505 14332 21539
rect 14280 21496 14332 21505
rect 14556 21496 14608 21548
rect 16580 21496 16632 21548
rect 17592 21496 17644 21548
rect 17960 21539 18012 21548
rect 17960 21505 17969 21539
rect 17969 21505 18003 21539
rect 18003 21505 18012 21539
rect 17960 21496 18012 21505
rect 18604 21564 18656 21616
rect 18788 21496 18840 21548
rect 18880 21496 18932 21548
rect 22376 21564 22428 21616
rect 30564 21632 30616 21684
rect 31484 21675 31536 21684
rect 31484 21641 31493 21675
rect 31493 21641 31527 21675
rect 31527 21641 31536 21675
rect 31484 21632 31536 21641
rect 31576 21632 31628 21684
rect 33416 21632 33468 21684
rect 35716 21675 35768 21684
rect 35716 21641 35725 21675
rect 35725 21641 35759 21675
rect 35759 21641 35768 21675
rect 35716 21632 35768 21641
rect 32036 21564 32088 21616
rect 35256 21564 35308 21616
rect 35808 21564 35860 21616
rect 25228 21496 25280 21548
rect 28816 21496 28868 21548
rect 29184 21539 29236 21548
rect 29184 21505 29193 21539
rect 29193 21505 29227 21539
rect 29227 21505 29236 21539
rect 29184 21496 29236 21505
rect 31116 21496 31168 21548
rect 15660 21428 15712 21480
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 17684 21428 17736 21480
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 15844 21360 15896 21412
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 19156 21428 19208 21480
rect 19340 21471 19392 21480
rect 19340 21437 19349 21471
rect 19349 21437 19383 21471
rect 19383 21437 19392 21471
rect 19340 21428 19392 21437
rect 20076 21428 20128 21480
rect 24400 21428 24452 21480
rect 24676 21471 24728 21480
rect 24676 21437 24685 21471
rect 24685 21437 24719 21471
rect 24719 21437 24728 21471
rect 24676 21428 24728 21437
rect 32680 21539 32732 21548
rect 32680 21505 32689 21539
rect 32689 21505 32723 21539
rect 32723 21505 32732 21539
rect 32680 21496 32732 21505
rect 32864 21539 32916 21548
rect 32864 21505 32873 21539
rect 32873 21505 32907 21539
rect 32907 21505 32916 21539
rect 32864 21496 32916 21505
rect 33692 21539 33744 21548
rect 33692 21505 33701 21539
rect 33701 21505 33735 21539
rect 33735 21505 33744 21539
rect 33692 21496 33744 21505
rect 34704 21496 34756 21548
rect 22376 21360 22428 21412
rect 16212 21292 16264 21344
rect 17408 21292 17460 21344
rect 18972 21292 19024 21344
rect 25964 21292 26016 21344
rect 26056 21335 26108 21344
rect 26056 21301 26065 21335
rect 26065 21301 26099 21335
rect 26099 21301 26108 21335
rect 26056 21292 26108 21301
rect 27252 21292 27304 21344
rect 28264 21292 28316 21344
rect 28816 21292 28868 21344
rect 32404 21428 32456 21480
rect 32588 21428 32640 21480
rect 35440 21539 35492 21548
rect 35440 21505 35449 21539
rect 35449 21505 35483 21539
rect 35483 21505 35492 21539
rect 35440 21496 35492 21505
rect 36176 21496 36228 21548
rect 38660 21496 38712 21548
rect 38844 21471 38896 21480
rect 38844 21437 38853 21471
rect 38853 21437 38887 21471
rect 38887 21437 38896 21471
rect 38844 21428 38896 21437
rect 31300 21403 31352 21412
rect 31300 21369 31309 21403
rect 31309 21369 31343 21403
rect 31343 21369 31352 21403
rect 31300 21360 31352 21369
rect 34796 21360 34848 21412
rect 35532 21360 35584 21412
rect 35808 21360 35860 21412
rect 38016 21360 38068 21412
rect 31852 21292 31904 21344
rect 33416 21292 33468 21344
rect 34428 21292 34480 21344
rect 34612 21292 34664 21344
rect 35440 21292 35492 21344
rect 38752 21292 38804 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7748 21131 7800 21140
rect 7748 21097 7757 21131
rect 7757 21097 7791 21131
rect 7791 21097 7800 21131
rect 7748 21088 7800 21097
rect 7840 21088 7892 21140
rect 14556 21088 14608 21140
rect 15660 21131 15712 21140
rect 15660 21097 15669 21131
rect 15669 21097 15703 21131
rect 15703 21097 15712 21131
rect 15660 21088 15712 21097
rect 16856 21088 16908 21140
rect 17592 21088 17644 21140
rect 18604 21088 18656 21140
rect 19340 21088 19392 21140
rect 25228 21131 25280 21140
rect 7656 21020 7708 21072
rect 9312 21020 9364 21072
rect 1492 20952 1544 21004
rect 2872 20952 2924 21004
rect 13360 20952 13412 21004
rect 15660 20952 15712 21004
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 19616 21020 19668 21072
rect 25228 21097 25237 21131
rect 25237 21097 25271 21131
rect 25271 21097 25280 21131
rect 25228 21088 25280 21097
rect 25964 21088 26016 21140
rect 38292 21131 38344 21140
rect 38292 21097 38301 21131
rect 38301 21097 38335 21131
rect 38335 21097 38344 21131
rect 38292 21088 38344 21097
rect 35808 21020 35860 21072
rect 19524 20995 19576 21004
rect 19524 20961 19533 20995
rect 19533 20961 19567 20995
rect 19567 20961 19576 20995
rect 19524 20952 19576 20961
rect 2228 20884 2280 20936
rect 7012 20884 7064 20936
rect 7748 20884 7800 20936
rect 7840 20927 7892 20936
rect 7840 20893 7849 20927
rect 7849 20893 7883 20927
rect 7883 20893 7892 20927
rect 10508 20927 10560 20936
rect 7840 20884 7892 20893
rect 7564 20816 7616 20868
rect 8024 20893 8033 20912
rect 8033 20893 8067 20912
rect 8067 20893 8076 20912
rect 8024 20860 8076 20893
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 15844 20927 15896 20936
rect 15844 20893 15853 20927
rect 15853 20893 15887 20927
rect 15887 20893 15896 20927
rect 15844 20884 15896 20893
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 17500 20927 17552 20936
rect 12440 20816 12492 20868
rect 13728 20816 13780 20868
rect 2964 20748 3016 20800
rect 6920 20748 6972 20800
rect 8668 20748 8720 20800
rect 10692 20748 10744 20800
rect 11060 20748 11112 20800
rect 15568 20748 15620 20800
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 18696 20884 18748 20936
rect 19294 20884 19346 20936
rect 19708 20927 19760 20936
rect 19708 20893 19718 20927
rect 19718 20893 19752 20927
rect 19752 20893 19760 20927
rect 19708 20884 19760 20893
rect 21640 20884 21692 20936
rect 28080 20952 28132 21004
rect 28264 20952 28316 21004
rect 32588 20995 32640 21004
rect 25780 20884 25832 20936
rect 26240 20884 26292 20936
rect 18144 20816 18196 20868
rect 19156 20816 19208 20868
rect 17868 20748 17920 20800
rect 22008 20816 22060 20868
rect 23020 20816 23072 20868
rect 26792 20816 26844 20868
rect 27252 20859 27304 20868
rect 27252 20825 27261 20859
rect 27261 20825 27295 20859
rect 27295 20825 27304 20859
rect 27252 20816 27304 20825
rect 27620 20884 27672 20936
rect 31576 20884 31628 20936
rect 32588 20961 32597 20995
rect 32597 20961 32631 20995
rect 32631 20961 32640 20995
rect 32588 20952 32640 20961
rect 32772 20952 32824 21004
rect 33600 20884 33652 20936
rect 34704 20884 34756 20936
rect 34244 20816 34296 20868
rect 22376 20748 22428 20800
rect 23388 20748 23440 20800
rect 26056 20748 26108 20800
rect 27528 20748 27580 20800
rect 27988 20791 28040 20800
rect 27988 20757 27997 20791
rect 27997 20757 28031 20791
rect 28031 20757 28040 20791
rect 27988 20748 28040 20757
rect 28080 20748 28132 20800
rect 34796 20748 34848 20800
rect 35348 20859 35400 20868
rect 35348 20825 35357 20859
rect 35357 20825 35391 20859
rect 35391 20825 35400 20859
rect 35348 20816 35400 20825
rect 35440 20859 35492 20868
rect 35440 20825 35449 20859
rect 35449 20825 35483 20859
rect 35483 20825 35492 20859
rect 35808 20884 35860 20936
rect 36268 20927 36320 20936
rect 36268 20893 36278 20927
rect 36278 20893 36312 20927
rect 36312 20893 36320 20927
rect 36268 20884 36320 20893
rect 35440 20816 35492 20825
rect 36360 20816 36412 20868
rect 36544 20859 36596 20868
rect 36544 20825 36553 20859
rect 36553 20825 36587 20859
rect 36587 20825 36596 20859
rect 36544 20816 36596 20825
rect 35808 20748 35860 20800
rect 36176 20748 36228 20800
rect 38752 20927 38804 20936
rect 38752 20893 38761 20927
rect 38761 20893 38795 20927
rect 38795 20893 38804 20927
rect 38752 20884 38804 20893
rect 37832 20816 37884 20868
rect 39856 20816 39908 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 2412 20544 2464 20596
rect 2964 20544 3016 20596
rect 8024 20544 8076 20596
rect 10508 20544 10560 20596
rect 11060 20544 11112 20596
rect 19294 20544 19346 20596
rect 8116 20476 8168 20528
rect 12440 20519 12492 20528
rect 12440 20485 12449 20519
rect 12449 20485 12483 20519
rect 12483 20485 12492 20519
rect 12900 20519 12952 20528
rect 12440 20476 12492 20485
rect 12900 20485 12909 20519
rect 12909 20485 12943 20519
rect 12943 20485 12952 20519
rect 12900 20476 12952 20485
rect 13176 20476 13228 20528
rect 16948 20476 17000 20528
rect 20168 20544 20220 20596
rect 22376 20587 22428 20596
rect 21732 20476 21784 20528
rect 22008 20519 22060 20528
rect 22008 20485 22017 20519
rect 22017 20485 22051 20519
rect 22051 20485 22060 20519
rect 22008 20476 22060 20485
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 25780 20587 25832 20596
rect 25780 20553 25789 20587
rect 25789 20553 25823 20587
rect 25823 20553 25832 20587
rect 25780 20544 25832 20553
rect 27620 20544 27672 20596
rect 27712 20544 27764 20596
rect 34060 20544 34112 20596
rect 3332 20408 3384 20460
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 7012 20451 7064 20460
rect 7012 20417 7021 20451
rect 7021 20417 7055 20451
rect 7055 20417 7064 20451
rect 7012 20408 7064 20417
rect 7840 20408 7892 20460
rect 8852 20408 8904 20460
rect 11796 20408 11848 20460
rect 16580 20408 16632 20460
rect 17132 20408 17184 20460
rect 2596 20383 2648 20392
rect 2596 20349 2605 20383
rect 2605 20349 2639 20383
rect 2639 20349 2648 20383
rect 2596 20340 2648 20349
rect 2688 20383 2740 20392
rect 2688 20349 2697 20383
rect 2697 20349 2731 20383
rect 2731 20349 2740 20383
rect 7748 20383 7800 20392
rect 2688 20340 2740 20349
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 10416 20340 10468 20392
rect 9680 20272 9732 20324
rect 9864 20272 9916 20324
rect 10600 20272 10652 20324
rect 15476 20340 15528 20392
rect 18052 20408 18104 20460
rect 19248 20408 19300 20460
rect 19340 20408 19392 20460
rect 17868 20340 17920 20392
rect 14832 20272 14884 20324
rect 15108 20272 15160 20324
rect 15568 20272 15620 20324
rect 17960 20272 18012 20324
rect 18420 20383 18472 20392
rect 18420 20349 18429 20383
rect 18429 20349 18463 20383
rect 18463 20349 18472 20383
rect 19524 20383 19576 20392
rect 18420 20340 18472 20349
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 19708 20383 19760 20392
rect 19708 20349 19718 20383
rect 19718 20349 19752 20383
rect 19752 20349 19760 20383
rect 19892 20383 19944 20392
rect 19708 20340 19760 20349
rect 19892 20349 19901 20383
rect 19901 20349 19935 20383
rect 19935 20349 19944 20383
rect 19892 20340 19944 20349
rect 20076 20340 20128 20392
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22468 20451 22520 20460
rect 22192 20408 22244 20417
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 26148 20408 26200 20460
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27988 20476 28040 20528
rect 35348 20476 35400 20528
rect 36360 20544 36412 20596
rect 36452 20476 36504 20528
rect 34796 20408 34848 20460
rect 35716 20451 35768 20460
rect 35716 20417 35725 20451
rect 35725 20417 35759 20451
rect 35759 20417 35768 20451
rect 35716 20408 35768 20417
rect 27712 20340 27764 20392
rect 27896 20340 27948 20392
rect 36176 20451 36228 20460
rect 36176 20417 36190 20451
rect 36190 20417 36224 20451
rect 36224 20417 36228 20451
rect 36176 20408 36228 20417
rect 38752 20408 38804 20460
rect 38200 20340 38252 20392
rect 39120 20383 39172 20392
rect 39120 20349 39129 20383
rect 39129 20349 39163 20383
rect 39163 20349 39172 20383
rect 39120 20340 39172 20349
rect 23388 20272 23440 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 3608 20247 3660 20256
rect 3608 20213 3617 20247
rect 3617 20213 3651 20247
rect 3651 20213 3660 20247
rect 3608 20204 3660 20213
rect 7656 20247 7708 20256
rect 7656 20213 7665 20247
rect 7665 20213 7699 20247
rect 7699 20213 7708 20247
rect 7656 20204 7708 20213
rect 9588 20204 9640 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 20352 20204 20404 20256
rect 21732 20204 21784 20256
rect 29552 20204 29604 20256
rect 40040 20204 40092 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2596 20000 2648 20052
rect 3424 20000 3476 20052
rect 8300 20000 8352 20052
rect 11796 20043 11848 20052
rect 11796 20009 11805 20043
rect 11805 20009 11839 20043
rect 11839 20009 11848 20043
rect 11796 20000 11848 20009
rect 12900 20000 12952 20052
rect 15936 20000 15988 20052
rect 17500 20000 17552 20052
rect 24124 20000 24176 20052
rect 27160 20000 27212 20052
rect 38752 20043 38804 20052
rect 1492 19864 1544 19916
rect 6828 19864 6880 19916
rect 2780 19796 2832 19848
rect 3608 19796 3660 19848
rect 7104 19796 7156 19848
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 2136 19728 2188 19780
rect 6920 19771 6972 19780
rect 6920 19737 6929 19771
rect 6929 19737 6963 19771
rect 6963 19737 6972 19771
rect 7932 19796 7984 19848
rect 8024 19771 8076 19780
rect 6920 19728 6972 19737
rect 8024 19737 8033 19771
rect 8033 19737 8067 19771
rect 8067 19737 8076 19771
rect 8024 19728 8076 19737
rect 8116 19728 8168 19780
rect 10232 19864 10284 19916
rect 13728 19864 13780 19916
rect 15568 19907 15620 19916
rect 15568 19873 15577 19907
rect 15577 19873 15611 19907
rect 15611 19873 15620 19907
rect 15568 19864 15620 19873
rect 23020 19932 23072 19984
rect 10692 19839 10744 19848
rect 10692 19805 10726 19839
rect 10726 19805 10744 19839
rect 10692 19796 10744 19805
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 13636 19796 13688 19848
rect 15384 19796 15436 19848
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 7012 19660 7064 19712
rect 7932 19660 7984 19712
rect 15108 19660 15160 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 15384 19660 15436 19712
rect 15568 19728 15620 19780
rect 15936 19796 15988 19848
rect 18420 19864 18472 19916
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 19800 19864 19852 19916
rect 20260 19864 20312 19916
rect 22192 19864 22244 19916
rect 22468 19864 22520 19916
rect 28908 19932 28960 19984
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 16120 19728 16172 19780
rect 20168 19728 20220 19780
rect 15844 19660 15896 19712
rect 21640 19796 21692 19848
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 29000 19864 29052 19916
rect 29736 19864 29788 19916
rect 28816 19839 28868 19848
rect 20352 19728 20404 19780
rect 22376 19728 22428 19780
rect 24676 19771 24728 19780
rect 24676 19737 24710 19771
rect 24710 19737 24728 19771
rect 24676 19728 24728 19737
rect 26240 19728 26292 19780
rect 27160 19728 27212 19780
rect 27528 19728 27580 19780
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 29552 19839 29604 19848
rect 29552 19805 29561 19839
rect 29561 19805 29595 19839
rect 29595 19805 29604 19839
rect 29552 19796 29604 19805
rect 30564 19796 30616 19848
rect 30748 19839 30800 19848
rect 30748 19805 30757 19839
rect 30757 19805 30791 19839
rect 30791 19805 30800 19839
rect 30748 19796 30800 19805
rect 38752 20009 38761 20043
rect 38761 20009 38795 20043
rect 38795 20009 38804 20043
rect 38752 20000 38804 20009
rect 39120 20000 39172 20052
rect 40500 20000 40552 20052
rect 31208 19907 31260 19916
rect 31208 19873 31217 19907
rect 31217 19873 31251 19907
rect 31251 19873 31260 19907
rect 31208 19864 31260 19873
rect 35808 19839 35860 19848
rect 25044 19660 25096 19712
rect 26148 19660 26200 19712
rect 29092 19660 29144 19712
rect 29736 19660 29788 19712
rect 30104 19660 30156 19712
rect 32588 19703 32640 19712
rect 32588 19669 32597 19703
rect 32597 19669 32631 19703
rect 32631 19669 32640 19703
rect 32588 19660 32640 19669
rect 35808 19805 35817 19839
rect 35817 19805 35851 19839
rect 35851 19805 35860 19839
rect 35808 19796 35860 19805
rect 36268 19839 36320 19848
rect 36268 19805 36282 19839
rect 36282 19805 36316 19839
rect 36316 19805 36320 19839
rect 38016 19839 38068 19848
rect 36268 19796 36320 19805
rect 38016 19805 38025 19839
rect 38025 19805 38059 19839
rect 38059 19805 38068 19839
rect 38016 19796 38068 19805
rect 38844 19864 38896 19916
rect 39120 19907 39172 19916
rect 39120 19873 39129 19907
rect 39129 19873 39163 19907
rect 39163 19873 39172 19907
rect 39120 19864 39172 19873
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 39028 19839 39080 19848
rect 39028 19805 39037 19839
rect 39037 19805 39071 19839
rect 39071 19805 39080 19839
rect 39028 19796 39080 19805
rect 34796 19728 34848 19780
rect 36084 19771 36136 19780
rect 36084 19737 36093 19771
rect 36093 19737 36127 19771
rect 36127 19737 36136 19771
rect 36084 19728 36136 19737
rect 37096 19728 37148 19780
rect 38200 19771 38252 19780
rect 38200 19737 38209 19771
rect 38209 19737 38243 19771
rect 38243 19737 38252 19771
rect 38200 19728 38252 19737
rect 39120 19660 39172 19712
rect 48320 19660 48372 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 5172 19388 5224 19440
rect 7840 19456 7892 19508
rect 1400 19320 1452 19372
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 3332 19320 3384 19372
rect 6920 19320 6972 19372
rect 7104 19320 7156 19372
rect 8208 19388 8260 19440
rect 8300 19320 8352 19372
rect 9404 19320 9456 19372
rect 11796 19388 11848 19440
rect 13544 19456 13596 19508
rect 15384 19456 15436 19508
rect 15936 19456 15988 19508
rect 17040 19456 17092 19508
rect 24676 19499 24728 19508
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 27344 19499 27396 19508
rect 16120 19388 16172 19440
rect 17408 19388 17460 19440
rect 27344 19465 27353 19499
rect 27353 19465 27387 19499
rect 27387 19465 27396 19499
rect 27344 19456 27396 19465
rect 30748 19456 30800 19508
rect 34060 19499 34112 19508
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 12348 19320 12400 19372
rect 12900 19320 12952 19372
rect 8116 19184 8168 19236
rect 13360 19320 13412 19372
rect 13636 19320 13688 19372
rect 15292 19363 15344 19372
rect 15292 19329 15301 19363
rect 15301 19329 15335 19363
rect 15335 19329 15344 19363
rect 15292 19320 15344 19329
rect 17132 19363 17184 19372
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 13452 19184 13504 19236
rect 2688 19116 2740 19168
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 7288 19116 7340 19168
rect 8024 19116 8076 19168
rect 16120 19252 16172 19304
rect 17132 19329 17141 19363
rect 17141 19329 17175 19363
rect 17175 19329 17184 19363
rect 17132 19320 17184 19329
rect 18328 19320 18380 19372
rect 19248 19320 19300 19372
rect 19156 19252 19208 19304
rect 19524 19252 19576 19304
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 21640 19320 21692 19372
rect 22100 19363 22152 19372
rect 22100 19329 22134 19363
rect 22134 19329 22152 19363
rect 22100 19320 22152 19329
rect 25136 19363 25188 19372
rect 25136 19329 25145 19363
rect 25145 19329 25179 19363
rect 25179 19329 25188 19363
rect 25136 19320 25188 19329
rect 26240 19431 26292 19440
rect 26240 19397 26265 19431
rect 26265 19397 26292 19431
rect 26240 19388 26292 19397
rect 27160 19431 27212 19440
rect 27160 19397 27185 19431
rect 27185 19397 27212 19431
rect 27160 19388 27212 19397
rect 28724 19388 28776 19440
rect 19892 19252 19944 19261
rect 20904 19252 20956 19304
rect 27988 19320 28040 19372
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 29644 19363 29696 19372
rect 29644 19329 29653 19363
rect 29653 19329 29687 19363
rect 29687 19329 29696 19363
rect 29644 19320 29696 19329
rect 30196 19363 30248 19372
rect 30196 19329 30205 19363
rect 30205 19329 30239 19363
rect 30239 19329 30248 19363
rect 30196 19320 30248 19329
rect 30656 19320 30708 19372
rect 28540 19252 28592 19304
rect 30472 19252 30524 19304
rect 30564 19252 30616 19304
rect 31116 19320 31168 19372
rect 32036 19320 32088 19372
rect 32588 19320 32640 19372
rect 34060 19465 34069 19499
rect 34069 19465 34103 19499
rect 34103 19465 34112 19499
rect 34060 19456 34112 19465
rect 39028 19456 39080 19508
rect 34152 19388 34204 19440
rect 31576 19295 31628 19304
rect 31576 19261 31585 19295
rect 31585 19261 31619 19295
rect 31619 19261 31628 19295
rect 31576 19252 31628 19261
rect 32220 19252 32272 19304
rect 15844 19184 15896 19236
rect 20812 19184 20864 19236
rect 25504 19184 25556 19236
rect 18052 19116 18104 19168
rect 18420 19116 18472 19168
rect 19892 19116 19944 19168
rect 20076 19116 20128 19168
rect 20996 19116 21048 19168
rect 22560 19116 22612 19168
rect 31944 19184 31996 19236
rect 32036 19184 32088 19236
rect 33876 19363 33928 19372
rect 33876 19329 33890 19363
rect 33890 19329 33924 19363
rect 33924 19329 33928 19363
rect 33876 19320 33928 19329
rect 35348 19320 35400 19372
rect 38292 19320 38344 19372
rect 40040 19388 40092 19440
rect 34796 19252 34848 19304
rect 38200 19252 38252 19304
rect 38016 19184 38068 19236
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 27068 19116 27120 19168
rect 29368 19116 29420 19168
rect 30012 19116 30064 19168
rect 36084 19116 36136 19168
rect 37004 19116 37056 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3148 18955 3200 18964
rect 3148 18921 3157 18955
rect 3157 18921 3191 18955
rect 3191 18921 3200 18955
rect 3148 18912 3200 18921
rect 7012 18912 7064 18964
rect 7380 18912 7432 18964
rect 17132 18912 17184 18964
rect 19524 18955 19576 18964
rect 19524 18921 19533 18955
rect 19533 18921 19567 18955
rect 19567 18921 19576 18955
rect 19524 18912 19576 18921
rect 1492 18708 1544 18760
rect 7748 18844 7800 18896
rect 6920 18776 6972 18828
rect 8852 18776 8904 18828
rect 7380 18708 7432 18760
rect 7932 18708 7984 18760
rect 8668 18708 8720 18760
rect 12532 18844 12584 18896
rect 15844 18844 15896 18896
rect 17040 18844 17092 18896
rect 17960 18844 18012 18896
rect 19892 18912 19944 18964
rect 20536 18955 20588 18964
rect 20536 18921 20545 18955
rect 20545 18921 20579 18955
rect 20579 18921 20588 18955
rect 20536 18912 20588 18921
rect 22100 18912 22152 18964
rect 22376 18912 22428 18964
rect 28724 18912 28776 18964
rect 28816 18955 28868 18964
rect 28816 18921 28825 18955
rect 28825 18921 28859 18955
rect 28859 18921 28868 18955
rect 29000 18955 29052 18964
rect 28816 18912 28868 18921
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 30196 18912 30248 18964
rect 30472 18912 30524 18964
rect 36636 18912 36688 18964
rect 25136 18844 25188 18896
rect 25412 18887 25464 18896
rect 25412 18853 25421 18887
rect 25421 18853 25455 18887
rect 25455 18853 25464 18887
rect 25412 18844 25464 18853
rect 28908 18844 28960 18896
rect 12532 18751 12584 18760
rect 3792 18640 3844 18692
rect 8208 18683 8260 18692
rect 8208 18649 8217 18683
rect 8217 18649 8251 18683
rect 8251 18649 8260 18683
rect 8208 18640 8260 18649
rect 10692 18640 10744 18692
rect 1768 18572 1820 18624
rect 6828 18572 6880 18624
rect 6920 18572 6972 18624
rect 10232 18572 10284 18624
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 18604 18776 18656 18828
rect 20260 18776 20312 18828
rect 22192 18776 22244 18828
rect 17316 18708 17368 18760
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 20720 18751 20772 18760
rect 15568 18683 15620 18692
rect 15568 18649 15577 18683
rect 15577 18649 15611 18683
rect 15611 18649 15620 18683
rect 15568 18640 15620 18649
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 12900 18572 12952 18624
rect 15752 18572 15804 18624
rect 15936 18572 15988 18624
rect 19248 18640 19300 18692
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 20996 18751 21048 18760
rect 20996 18717 21005 18751
rect 21005 18717 21039 18751
rect 21039 18717 21048 18751
rect 20996 18708 21048 18717
rect 22560 18776 22612 18828
rect 30104 18776 30156 18828
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22652 18751 22704 18760
rect 22376 18708 22428 18717
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 25136 18640 25188 18692
rect 26148 18640 26200 18692
rect 28632 18683 28684 18692
rect 28632 18649 28641 18683
rect 28641 18649 28675 18683
rect 28675 18649 28684 18683
rect 28632 18640 28684 18649
rect 29184 18708 29236 18760
rect 30012 18751 30064 18760
rect 31852 18776 31904 18828
rect 30012 18717 30026 18751
rect 30026 18717 30060 18751
rect 30060 18717 30064 18751
rect 30012 18708 30064 18717
rect 30932 18708 30984 18760
rect 32036 18751 32088 18760
rect 32036 18717 32045 18751
rect 32045 18717 32079 18751
rect 32079 18717 32088 18751
rect 32036 18708 32088 18717
rect 32220 18751 32272 18760
rect 32220 18717 32227 18751
rect 32227 18717 32272 18751
rect 32220 18708 32272 18717
rect 33508 18776 33560 18828
rect 36176 18844 36228 18896
rect 38660 18844 38712 18896
rect 32772 18708 32824 18760
rect 33876 18708 33928 18760
rect 35992 18751 36044 18760
rect 35992 18717 36001 18751
rect 36001 18717 36035 18751
rect 36035 18717 36044 18751
rect 35992 18708 36044 18717
rect 36636 18708 36688 18760
rect 37188 18751 37240 18760
rect 37188 18717 37197 18751
rect 37197 18717 37231 18751
rect 37231 18717 37240 18751
rect 37188 18708 37240 18717
rect 37372 18751 37424 18760
rect 37372 18717 37379 18751
rect 37379 18717 37424 18751
rect 37372 18708 37424 18717
rect 40040 18751 40092 18760
rect 40040 18717 40049 18751
rect 40049 18717 40083 18751
rect 40083 18717 40092 18751
rect 40040 18708 40092 18717
rect 29552 18640 29604 18692
rect 22560 18615 22612 18624
rect 22560 18581 22569 18615
rect 22569 18581 22603 18615
rect 22603 18581 22612 18615
rect 22560 18572 22612 18581
rect 24400 18572 24452 18624
rect 27068 18572 27120 18624
rect 27896 18572 27948 18624
rect 29460 18572 29512 18624
rect 36912 18640 36964 18692
rect 37004 18640 37056 18692
rect 37556 18683 37608 18692
rect 37556 18649 37565 18683
rect 37565 18649 37599 18683
rect 37599 18649 37608 18683
rect 37556 18640 37608 18649
rect 39948 18640 40000 18692
rect 32588 18572 32640 18624
rect 36084 18572 36136 18624
rect 36636 18615 36688 18624
rect 36636 18581 36645 18615
rect 36645 18581 36679 18615
rect 36679 18581 36688 18615
rect 36636 18572 36688 18581
rect 37832 18615 37884 18624
rect 37832 18581 37841 18615
rect 37841 18581 37875 18615
rect 37875 18581 37884 18615
rect 37832 18572 37884 18581
rect 38016 18572 38068 18624
rect 40408 18615 40460 18624
rect 40408 18581 40417 18615
rect 40417 18581 40451 18615
rect 40451 18581 40460 18615
rect 40408 18572 40460 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 3148 18368 3200 18420
rect 3884 18411 3936 18420
rect 3884 18377 3893 18411
rect 3893 18377 3927 18411
rect 3927 18377 3936 18411
rect 3884 18368 3936 18377
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 15568 18368 15620 18420
rect 17224 18368 17276 18420
rect 18328 18368 18380 18420
rect 20720 18368 20772 18420
rect 20812 18368 20864 18420
rect 37832 18368 37884 18420
rect 2688 18343 2740 18352
rect 2688 18309 2697 18343
rect 2697 18309 2731 18343
rect 2731 18309 2740 18343
rect 2688 18300 2740 18309
rect 4620 18232 4672 18284
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7840 18232 7892 18284
rect 10140 18300 10192 18352
rect 15752 18300 15804 18352
rect 8944 18232 8996 18284
rect 12348 18232 12400 18284
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 16120 18232 16172 18284
rect 16672 18232 16724 18284
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18604 18232 18656 18284
rect 19064 18232 19116 18284
rect 3056 18164 3108 18216
rect 3884 18164 3936 18216
rect 11428 18164 11480 18216
rect 15200 18164 15252 18216
rect 6184 18096 6236 18148
rect 14464 18096 14516 18148
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 17960 18164 18012 18216
rect 3332 18028 3384 18080
rect 8024 18028 8076 18080
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 19248 18207 19300 18216
rect 18144 18164 18196 18173
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 22376 18300 22428 18352
rect 19984 18232 20036 18284
rect 22008 18232 22060 18284
rect 20444 18207 20496 18216
rect 19064 18096 19116 18148
rect 20444 18173 20453 18207
rect 20453 18173 20487 18207
rect 20487 18173 20496 18207
rect 20444 18164 20496 18173
rect 20628 18164 20680 18216
rect 30840 18300 30892 18352
rect 31208 18343 31260 18352
rect 31208 18309 31217 18343
rect 31217 18309 31251 18343
rect 31251 18309 31260 18343
rect 31208 18300 31260 18309
rect 31576 18300 31628 18352
rect 37372 18300 37424 18352
rect 27068 18275 27120 18284
rect 27068 18241 27077 18275
rect 27077 18241 27111 18275
rect 27111 18241 27120 18275
rect 27068 18232 27120 18241
rect 27160 18232 27212 18284
rect 29184 18275 29236 18284
rect 18144 18028 18196 18080
rect 18328 18028 18380 18080
rect 21548 18028 21600 18080
rect 22284 18096 22336 18148
rect 28632 18164 28684 18216
rect 29184 18241 29193 18275
rect 29193 18241 29227 18275
rect 29227 18241 29236 18275
rect 29184 18232 29236 18241
rect 29460 18232 29512 18284
rect 30380 18232 30432 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 31116 18275 31168 18284
rect 31116 18241 31123 18275
rect 31123 18241 31168 18275
rect 31116 18232 31168 18241
rect 31668 18232 31720 18284
rect 33508 18232 33560 18284
rect 35808 18232 35860 18284
rect 35992 18232 36044 18284
rect 37188 18232 37240 18284
rect 32128 18164 32180 18216
rect 33876 18207 33928 18216
rect 22192 18028 22244 18080
rect 30288 18096 30340 18148
rect 30380 18096 30432 18148
rect 33876 18173 33885 18207
rect 33885 18173 33919 18207
rect 33919 18173 33928 18207
rect 33876 18164 33928 18173
rect 34796 18164 34848 18216
rect 37464 18275 37516 18284
rect 37464 18241 37473 18275
rect 37473 18241 37507 18275
rect 37507 18241 37516 18275
rect 38936 18300 38988 18352
rect 39948 18300 40000 18352
rect 37464 18232 37516 18241
rect 38016 18164 38068 18216
rect 38200 18164 38252 18216
rect 33968 18096 34020 18148
rect 40040 18232 40092 18284
rect 40408 18164 40460 18216
rect 40500 18207 40552 18216
rect 40500 18173 40509 18207
rect 40509 18173 40543 18207
rect 40543 18173 40552 18207
rect 40500 18164 40552 18173
rect 29552 18028 29604 18080
rect 31484 18028 31536 18080
rect 37372 18071 37424 18080
rect 37372 18037 37381 18071
rect 37381 18037 37415 18071
rect 37415 18037 37424 18071
rect 37372 18028 37424 18037
rect 40316 18028 40368 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 6184 17867 6236 17876
rect 3792 17799 3844 17808
rect 3792 17765 3801 17799
rect 3801 17765 3835 17799
rect 3835 17765 3844 17799
rect 3792 17756 3844 17765
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 8944 17867 8996 17876
rect 8944 17833 8953 17867
rect 8953 17833 8987 17867
rect 8987 17833 8996 17867
rect 8944 17824 8996 17833
rect 12624 17756 12676 17808
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 3332 17620 3384 17672
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 9496 17688 9548 17740
rect 15660 17824 15712 17876
rect 16212 17824 16264 17876
rect 18236 17824 18288 17876
rect 26240 17824 26292 17876
rect 27160 17867 27212 17876
rect 27160 17833 27169 17867
rect 27169 17833 27203 17867
rect 27203 17833 27212 17867
rect 27160 17824 27212 17833
rect 29000 17824 29052 17876
rect 30288 17824 30340 17876
rect 31484 17824 31536 17876
rect 21548 17756 21600 17808
rect 18512 17731 18564 17740
rect 9128 17663 9180 17672
rect 6736 17552 6788 17604
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 9220 17620 9272 17672
rect 9680 17620 9732 17672
rect 12256 17620 12308 17672
rect 12716 17620 12768 17672
rect 13360 17620 13412 17672
rect 13820 17620 13872 17672
rect 18512 17697 18521 17731
rect 18521 17697 18555 17731
rect 18555 17697 18564 17731
rect 18512 17688 18564 17697
rect 18788 17688 18840 17740
rect 23940 17688 23992 17740
rect 24400 17731 24452 17740
rect 24400 17697 24409 17731
rect 24409 17697 24443 17731
rect 24443 17697 24452 17731
rect 24400 17688 24452 17697
rect 32036 17756 32088 17808
rect 27436 17688 27488 17740
rect 31208 17688 31260 17740
rect 31852 17688 31904 17740
rect 16120 17620 16172 17672
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18420 17620 18472 17629
rect 18696 17620 18748 17672
rect 19984 17620 20036 17672
rect 21640 17663 21692 17672
rect 21640 17629 21649 17663
rect 21649 17629 21683 17663
rect 21683 17629 21692 17663
rect 21640 17620 21692 17629
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 12992 17595 13044 17604
rect 9312 17552 9364 17561
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 6184 17484 6236 17536
rect 7472 17484 7524 17536
rect 9128 17484 9180 17536
rect 9496 17484 9548 17536
rect 12164 17484 12216 17536
rect 12992 17561 13001 17595
rect 13001 17561 13035 17595
rect 13035 17561 13044 17595
rect 12992 17552 13044 17561
rect 15292 17552 15344 17604
rect 17132 17552 17184 17604
rect 14740 17484 14792 17536
rect 15108 17484 15160 17536
rect 18144 17484 18196 17536
rect 21916 17595 21968 17604
rect 21916 17561 21950 17595
rect 21950 17561 21968 17595
rect 21916 17552 21968 17561
rect 24676 17595 24728 17604
rect 24676 17561 24710 17595
rect 24710 17561 24728 17595
rect 27068 17663 27120 17672
rect 27068 17629 27077 17663
rect 27077 17629 27111 17663
rect 27111 17629 27120 17663
rect 29552 17663 29604 17672
rect 27068 17620 27120 17629
rect 29552 17629 29561 17663
rect 29561 17629 29595 17663
rect 29595 17629 29604 17663
rect 29552 17620 29604 17629
rect 30564 17620 30616 17672
rect 32404 17620 32456 17672
rect 34796 17620 34848 17672
rect 37464 17824 37516 17876
rect 40040 17824 40092 17876
rect 48320 17867 48372 17876
rect 38016 17688 38068 17740
rect 40500 17688 40552 17740
rect 41052 17688 41104 17740
rect 48320 17833 48329 17867
rect 48329 17833 48363 17867
rect 48363 17833 48372 17867
rect 48320 17824 48372 17833
rect 48596 17824 48648 17876
rect 37372 17663 37424 17672
rect 37372 17629 37381 17663
rect 37381 17629 37415 17663
rect 37415 17629 37424 17663
rect 37372 17620 37424 17629
rect 40040 17663 40092 17672
rect 24676 17552 24728 17561
rect 33692 17552 33744 17604
rect 34060 17552 34112 17604
rect 40040 17629 40049 17663
rect 40049 17629 40083 17663
rect 40083 17629 40092 17663
rect 40040 17620 40092 17629
rect 40316 17663 40368 17672
rect 40316 17629 40325 17663
rect 40325 17629 40359 17663
rect 40359 17629 40368 17663
rect 40316 17620 40368 17629
rect 42892 17595 42944 17604
rect 42892 17561 42926 17595
rect 42926 17561 42944 17595
rect 42892 17552 42944 17561
rect 20628 17484 20680 17536
rect 22376 17484 22428 17536
rect 25228 17484 25280 17536
rect 34704 17484 34756 17536
rect 35992 17484 36044 17536
rect 37188 17484 37240 17536
rect 39856 17484 39908 17536
rect 43996 17527 44048 17536
rect 43996 17493 44005 17527
rect 44005 17493 44039 17527
rect 44039 17493 44048 17527
rect 43996 17484 44048 17493
rect 45284 17552 45336 17604
rect 47860 17552 47912 17604
rect 47124 17484 47176 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 6828 17280 6880 17332
rect 15108 17280 15160 17332
rect 15292 17323 15344 17332
rect 15292 17289 15301 17323
rect 15301 17289 15335 17323
rect 15335 17289 15344 17323
rect 15292 17280 15344 17289
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 16120 17280 16172 17332
rect 22192 17280 22244 17332
rect 22376 17323 22428 17332
rect 22376 17289 22385 17323
rect 22385 17289 22419 17323
rect 22419 17289 22428 17323
rect 22376 17280 22428 17289
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 1952 17212 2004 17264
rect 2412 17144 2464 17196
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 18420 17212 18472 17264
rect 25504 17280 25556 17332
rect 27068 17280 27120 17332
rect 30288 17280 30340 17332
rect 32680 17280 32732 17332
rect 38936 17323 38988 17332
rect 38936 17289 38945 17323
rect 38945 17289 38979 17323
rect 38979 17289 38988 17323
rect 38936 17280 38988 17289
rect 42892 17323 42944 17332
rect 42892 17289 42901 17323
rect 42901 17289 42935 17323
rect 42935 17289 42944 17323
rect 42892 17280 42944 17289
rect 45284 17323 45336 17332
rect 45284 17289 45293 17323
rect 45293 17289 45327 17323
rect 45327 17289 45336 17323
rect 45284 17280 45336 17289
rect 7840 17144 7892 17196
rect 8944 17144 8996 17196
rect 9128 17144 9180 17196
rect 10140 17144 10192 17196
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 6644 17076 6696 17128
rect 15384 17144 15436 17196
rect 18512 17144 18564 17196
rect 19064 17144 19116 17196
rect 19156 17144 19208 17196
rect 22284 17144 22336 17196
rect 22652 17144 22704 17196
rect 28908 17212 28960 17264
rect 31852 17212 31904 17264
rect 26056 17187 26108 17196
rect 26056 17153 26065 17187
rect 26065 17153 26099 17187
rect 26099 17153 26108 17187
rect 26056 17144 26108 17153
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 26884 17144 26936 17196
rect 27436 17187 27488 17196
rect 27436 17153 27445 17187
rect 27445 17153 27479 17187
rect 27479 17153 27488 17187
rect 27436 17144 27488 17153
rect 27528 17144 27580 17196
rect 29828 17144 29880 17196
rect 30932 17187 30984 17196
rect 30932 17153 30941 17187
rect 30941 17153 30975 17187
rect 30975 17153 30984 17187
rect 30932 17144 30984 17153
rect 31116 17187 31168 17196
rect 31116 17153 31123 17187
rect 31123 17153 31168 17187
rect 31116 17144 31168 17153
rect 31300 17187 31352 17196
rect 31300 17153 31309 17187
rect 31309 17153 31343 17187
rect 31343 17153 31352 17187
rect 31300 17144 31352 17153
rect 17132 17076 17184 17128
rect 17500 17076 17552 17128
rect 18604 17076 18656 17128
rect 21916 17076 21968 17128
rect 22100 17076 22152 17128
rect 1676 17008 1728 17060
rect 1400 16940 1452 16992
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 7472 16940 7524 16992
rect 11980 17008 12032 17060
rect 12256 17008 12308 17060
rect 24676 17008 24728 17060
rect 25044 17076 25096 17128
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 25504 17076 25556 17128
rect 30288 17076 30340 17128
rect 32036 17144 32088 17196
rect 32220 17187 32272 17196
rect 32220 17153 32230 17187
rect 32230 17153 32264 17187
rect 32264 17153 32272 17187
rect 32220 17144 32272 17153
rect 31668 17076 31720 17128
rect 32772 17144 32824 17196
rect 37280 17144 37332 17196
rect 43076 17187 43128 17196
rect 43076 17153 43085 17187
rect 43085 17153 43119 17187
rect 43119 17153 43128 17187
rect 43076 17144 43128 17153
rect 45560 17144 45612 17196
rect 37372 17076 37424 17128
rect 25688 17008 25740 17060
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 12716 16940 12768 16992
rect 13912 16940 13964 16992
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 15384 16940 15436 16992
rect 40040 16940 40092 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2044 16736 2096 16788
rect 8944 16779 8996 16788
rect 8944 16745 8953 16779
rect 8953 16745 8987 16779
rect 8987 16745 8996 16779
rect 8944 16736 8996 16745
rect 12256 16779 12308 16788
rect 1492 16532 1544 16584
rect 1952 16532 2004 16584
rect 2504 16532 2556 16584
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 2780 16396 2832 16448
rect 4896 16464 4948 16516
rect 8116 16464 8168 16516
rect 3792 16439 3844 16448
rect 3792 16405 3801 16439
rect 3801 16405 3835 16439
rect 3835 16405 3844 16439
rect 3792 16396 3844 16405
rect 6736 16396 6788 16448
rect 9220 16600 9272 16652
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 12256 16745 12265 16779
rect 12265 16745 12299 16779
rect 12299 16745 12308 16779
rect 12256 16736 12308 16745
rect 14648 16779 14700 16788
rect 14648 16745 14657 16779
rect 14657 16745 14691 16779
rect 14691 16745 14700 16779
rect 14648 16736 14700 16745
rect 14740 16736 14792 16788
rect 17040 16736 17092 16788
rect 11980 16668 12032 16720
rect 12992 16668 13044 16720
rect 13360 16711 13412 16720
rect 13360 16677 13369 16711
rect 13369 16677 13403 16711
rect 13403 16677 13412 16711
rect 13360 16668 13412 16677
rect 35624 16736 35676 16788
rect 43076 16779 43128 16788
rect 18880 16668 18932 16720
rect 22100 16668 22152 16720
rect 24676 16668 24728 16720
rect 27436 16668 27488 16720
rect 29368 16668 29420 16720
rect 31852 16668 31904 16720
rect 32864 16668 32916 16720
rect 43076 16745 43085 16779
rect 43085 16745 43119 16779
rect 43119 16745 43128 16779
rect 43076 16736 43128 16745
rect 45560 16779 45612 16788
rect 45560 16745 45569 16779
rect 45569 16745 45603 16779
rect 45603 16745 45612 16779
rect 45560 16736 45612 16745
rect 18328 16575 18380 16584
rect 18328 16541 18337 16575
rect 18337 16541 18371 16575
rect 18371 16541 18380 16575
rect 18328 16532 18380 16541
rect 18696 16532 18748 16584
rect 22192 16600 22244 16652
rect 24124 16532 24176 16584
rect 26056 16600 26108 16652
rect 37004 16643 37056 16652
rect 37004 16609 37013 16643
rect 37013 16609 37047 16643
rect 37047 16609 37056 16643
rect 37188 16643 37240 16652
rect 37004 16600 37056 16609
rect 37188 16609 37197 16643
rect 37197 16609 37231 16643
rect 37231 16609 37240 16643
rect 37188 16600 37240 16609
rect 24860 16532 24912 16584
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 26148 16532 26200 16584
rect 26516 16532 26568 16584
rect 9128 16396 9180 16448
rect 10784 16464 10836 16516
rect 13084 16464 13136 16516
rect 14556 16507 14608 16516
rect 14556 16473 14565 16507
rect 14565 16473 14599 16507
rect 14599 16473 14608 16507
rect 14556 16464 14608 16473
rect 15384 16464 15436 16516
rect 10876 16396 10928 16448
rect 12624 16396 12676 16448
rect 18420 16464 18472 16516
rect 29368 16464 29420 16516
rect 29552 16507 29604 16516
rect 29552 16473 29561 16507
rect 29561 16473 29595 16507
rect 29595 16473 29604 16507
rect 29552 16464 29604 16473
rect 29828 16464 29880 16516
rect 30380 16532 30432 16584
rect 30932 16575 30984 16584
rect 30932 16541 30941 16575
rect 30941 16541 30975 16575
rect 30975 16541 30984 16575
rect 30932 16532 30984 16541
rect 33784 16575 33836 16584
rect 33784 16541 33793 16575
rect 33793 16541 33827 16575
rect 33827 16541 33836 16575
rect 33784 16532 33836 16541
rect 33968 16575 34020 16584
rect 33968 16541 33977 16575
rect 33977 16541 34011 16575
rect 34011 16541 34020 16575
rect 33968 16532 34020 16541
rect 31208 16464 31260 16516
rect 34796 16464 34848 16516
rect 35992 16464 36044 16516
rect 37372 16600 37424 16652
rect 40224 16600 40276 16652
rect 43260 16600 43312 16652
rect 43996 16643 44048 16652
rect 43996 16609 44005 16643
rect 44005 16609 44039 16643
rect 44039 16609 44048 16643
rect 43996 16600 44048 16609
rect 40592 16532 40644 16584
rect 43720 16575 43772 16584
rect 43720 16541 43729 16575
rect 43729 16541 43763 16575
rect 43763 16541 43772 16575
rect 43720 16532 43772 16541
rect 43812 16575 43864 16584
rect 43812 16541 43821 16575
rect 43821 16541 43855 16575
rect 43855 16541 43864 16575
rect 45008 16643 45060 16652
rect 45008 16609 45017 16643
rect 45017 16609 45051 16643
rect 45051 16609 45060 16643
rect 45008 16600 45060 16609
rect 45468 16600 45520 16652
rect 43812 16532 43864 16541
rect 46572 16575 46624 16584
rect 46572 16541 46581 16575
rect 46581 16541 46615 16575
rect 46615 16541 46624 16575
rect 46572 16532 46624 16541
rect 40316 16507 40368 16516
rect 40316 16473 40325 16507
rect 40325 16473 40359 16507
rect 40359 16473 40368 16507
rect 40316 16464 40368 16473
rect 41236 16464 41288 16516
rect 45008 16464 45060 16516
rect 45100 16464 45152 16516
rect 22100 16396 22152 16448
rect 25320 16439 25372 16448
rect 25320 16405 25329 16439
rect 25329 16405 25363 16439
rect 25363 16405 25372 16439
rect 25320 16396 25372 16405
rect 29000 16396 29052 16448
rect 30748 16396 30800 16448
rect 33876 16439 33928 16448
rect 33876 16405 33885 16439
rect 33885 16405 33919 16439
rect 33919 16405 33928 16439
rect 33876 16396 33928 16405
rect 35532 16396 35584 16448
rect 37280 16396 37332 16448
rect 40960 16439 41012 16448
rect 40960 16405 40969 16439
rect 40969 16405 41003 16439
rect 41003 16405 41012 16439
rect 40960 16396 41012 16405
rect 45284 16439 45336 16448
rect 45284 16405 45293 16439
rect 45293 16405 45327 16439
rect 45327 16405 45336 16439
rect 45284 16396 45336 16405
rect 45468 16464 45520 16516
rect 47032 16507 47084 16516
rect 47032 16473 47066 16507
rect 47066 16473 47084 16507
rect 47032 16464 47084 16473
rect 47952 16439 48004 16448
rect 47952 16405 47961 16439
rect 47961 16405 47995 16439
rect 47995 16405 48004 16439
rect 47952 16396 48004 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2412 16235 2464 16244
rect 2412 16201 2421 16235
rect 2421 16201 2455 16235
rect 2455 16201 2464 16235
rect 2412 16192 2464 16201
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 2780 16192 2832 16201
rect 6644 16192 6696 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 10876 16192 10928 16244
rect 18328 16192 18380 16244
rect 2320 16124 2372 16176
rect 15384 16124 15436 16176
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 3792 16056 3844 16108
rect 6276 16056 6328 16108
rect 10508 16056 10560 16108
rect 14464 16056 14516 16108
rect 14924 16056 14976 16108
rect 18788 16124 18840 16176
rect 20904 16167 20956 16176
rect 20904 16133 20913 16167
rect 20913 16133 20947 16167
rect 20947 16133 20956 16167
rect 20904 16124 20956 16133
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 18236 16099 18288 16108
rect 17500 16056 17552 16065
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 18696 16056 18748 16108
rect 19064 16056 19116 16108
rect 24952 16192 25004 16244
rect 21640 16124 21692 16176
rect 24124 16124 24176 16176
rect 31116 16192 31168 16244
rect 21916 16056 21968 16108
rect 23940 16099 23992 16108
rect 23940 16065 23949 16099
rect 23949 16065 23983 16099
rect 23983 16065 23992 16099
rect 23940 16056 23992 16065
rect 24584 16056 24636 16108
rect 30472 16124 30524 16176
rect 33140 16235 33192 16244
rect 33140 16201 33149 16235
rect 33149 16201 33183 16235
rect 33183 16201 33192 16235
rect 33140 16192 33192 16201
rect 32128 16124 32180 16176
rect 28632 16056 28684 16108
rect 29000 16056 29052 16108
rect 29368 16056 29420 16108
rect 31116 16099 31168 16108
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 4804 15988 4856 16040
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 8116 15988 8168 16040
rect 11888 15988 11940 16040
rect 13820 15988 13872 16040
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 15752 15963 15804 15972
rect 15752 15929 15761 15963
rect 15761 15929 15795 15963
rect 15795 15929 15804 15963
rect 15752 15920 15804 15929
rect 17316 16031 17368 16040
rect 17316 15997 17325 16031
rect 17325 15997 17359 16031
rect 17359 15997 17368 16031
rect 17316 15988 17368 15997
rect 18788 15988 18840 16040
rect 18972 15988 19024 16040
rect 29276 16031 29328 16040
rect 19156 15920 19208 15972
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 31116 16065 31125 16099
rect 31125 16065 31159 16099
rect 31159 16065 31168 16099
rect 31116 16056 31168 16065
rect 32404 16056 32456 16108
rect 41144 16192 41196 16244
rect 45284 16192 45336 16244
rect 47032 16192 47084 16244
rect 34428 16167 34480 16176
rect 34428 16133 34462 16167
rect 34462 16133 34480 16167
rect 34428 16124 34480 16133
rect 34520 16124 34572 16176
rect 40960 16124 41012 16176
rect 43812 16124 43864 16176
rect 33876 16056 33928 16108
rect 40224 16056 40276 16108
rect 41052 16056 41104 16108
rect 43720 16056 43772 16108
rect 33324 16031 33376 16040
rect 33324 15997 33333 16031
rect 33333 15997 33367 16031
rect 33367 15997 33376 16031
rect 33324 15988 33376 15997
rect 26332 15920 26384 15972
rect 27988 15920 28040 15972
rect 7840 15852 7892 15904
rect 7932 15852 7984 15904
rect 8116 15852 8168 15904
rect 10876 15852 10928 15904
rect 18052 15852 18104 15904
rect 18972 15852 19024 15904
rect 19248 15852 19300 15904
rect 20352 15895 20404 15904
rect 20352 15861 20361 15895
rect 20361 15861 20395 15895
rect 20395 15861 20404 15895
rect 20352 15852 20404 15861
rect 22008 15852 22060 15904
rect 22192 15852 22244 15904
rect 26424 15852 26476 15904
rect 30288 15852 30340 15904
rect 30932 15852 30984 15904
rect 32128 15963 32180 15972
rect 32128 15929 32137 15963
rect 32137 15929 32171 15963
rect 32171 15929 32180 15963
rect 33968 15988 34020 16040
rect 45192 16056 45244 16108
rect 47952 16124 48004 16176
rect 46940 16056 46992 16108
rect 47584 16099 47636 16108
rect 47584 16065 47593 16099
rect 47593 16065 47627 16099
rect 47627 16065 47636 16099
rect 47584 16056 47636 16065
rect 48412 16056 48464 16108
rect 32128 15920 32180 15929
rect 46572 15920 46624 15972
rect 33508 15852 33560 15904
rect 41696 15895 41748 15904
rect 41696 15861 41705 15895
rect 41705 15861 41739 15895
rect 41739 15861 41748 15895
rect 41696 15852 41748 15861
rect 41972 15852 42024 15904
rect 45100 15852 45152 15904
rect 45192 15852 45244 15904
rect 47124 15852 47176 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15648 2188 15700
rect 6276 15691 6328 15700
rect 2872 15580 2924 15632
rect 3056 15512 3108 15564
rect 3516 15444 3568 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 5632 15376 5684 15428
rect 6276 15657 6285 15691
rect 6285 15657 6319 15691
rect 6319 15657 6328 15691
rect 6276 15648 6328 15657
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 14924 15691 14976 15700
rect 14924 15657 14933 15691
rect 14933 15657 14967 15691
rect 14967 15657 14976 15691
rect 14924 15648 14976 15657
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 17960 15648 18012 15700
rect 18236 15648 18288 15700
rect 18328 15648 18380 15700
rect 19064 15648 19116 15700
rect 19156 15648 19208 15700
rect 10600 15512 10652 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 18788 15580 18840 15632
rect 24124 15648 24176 15700
rect 24584 15691 24636 15700
rect 24584 15657 24593 15691
rect 24593 15657 24627 15691
rect 24627 15657 24636 15691
rect 24584 15648 24636 15657
rect 20260 15580 20312 15632
rect 26424 15648 26476 15700
rect 26608 15648 26660 15700
rect 18052 15512 18104 15564
rect 18604 15555 18656 15564
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 19064 15512 19116 15564
rect 6644 15487 6696 15496
rect 6644 15453 6653 15487
rect 6653 15453 6687 15487
rect 6687 15453 6696 15487
rect 6644 15444 6696 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 10876 15487 10928 15496
rect 6736 15444 6788 15453
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 18328 15487 18380 15496
rect 18328 15453 18337 15487
rect 18337 15453 18371 15487
rect 18371 15453 18380 15487
rect 18328 15444 18380 15453
rect 18512 15487 18564 15496
rect 18512 15453 18521 15487
rect 18521 15453 18555 15487
rect 18555 15453 18564 15487
rect 18512 15444 18564 15453
rect 18972 15444 19024 15496
rect 22008 15487 22060 15496
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 11060 15308 11112 15360
rect 15384 15376 15436 15428
rect 15752 15376 15804 15428
rect 16304 15308 16356 15360
rect 18604 15376 18656 15428
rect 19248 15376 19300 15428
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22192 15487 22244 15496
rect 22008 15444 22060 15453
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22652 15444 22704 15496
rect 24860 15512 24912 15564
rect 26608 15512 26660 15564
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 25412 15444 25464 15496
rect 29552 15648 29604 15700
rect 30748 15580 30800 15632
rect 33784 15648 33836 15700
rect 33968 15648 34020 15700
rect 40592 15691 40644 15700
rect 32772 15580 32824 15632
rect 21916 15376 21968 15428
rect 20352 15308 20404 15360
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 26516 15419 26568 15428
rect 26516 15385 26541 15419
rect 26541 15385 26568 15419
rect 26516 15376 26568 15385
rect 30196 15444 30248 15496
rect 30288 15487 30340 15496
rect 30288 15453 30297 15487
rect 30297 15453 30331 15487
rect 30331 15453 30340 15487
rect 30288 15444 30340 15453
rect 30564 15444 30616 15496
rect 32128 15444 32180 15496
rect 33508 15487 33560 15496
rect 33508 15453 33517 15487
rect 33517 15453 33551 15487
rect 33551 15453 33560 15487
rect 33508 15444 33560 15453
rect 34060 15512 34112 15564
rect 36268 15580 36320 15632
rect 37372 15580 37424 15632
rect 34796 15444 34848 15496
rect 27160 15419 27212 15428
rect 27160 15385 27169 15419
rect 27169 15385 27203 15419
rect 27203 15385 27212 15419
rect 27160 15376 27212 15385
rect 28264 15308 28316 15360
rect 30380 15376 30432 15428
rect 31300 15376 31352 15428
rect 31484 15376 31536 15428
rect 31024 15308 31076 15360
rect 31208 15308 31260 15360
rect 38660 15512 38712 15564
rect 40592 15657 40601 15691
rect 40601 15657 40635 15691
rect 40635 15657 40644 15691
rect 40592 15648 40644 15657
rect 54760 15691 54812 15700
rect 54760 15657 54769 15691
rect 54769 15657 54803 15691
rect 54803 15657 54812 15691
rect 54760 15648 54812 15657
rect 41696 15580 41748 15632
rect 35992 15487 36044 15496
rect 35992 15453 36001 15487
rect 36001 15453 36035 15487
rect 36035 15453 36044 15487
rect 35992 15444 36044 15453
rect 37924 15487 37976 15496
rect 37924 15453 37933 15487
rect 37933 15453 37967 15487
rect 37967 15453 37976 15487
rect 37924 15444 37976 15453
rect 41972 15555 42024 15564
rect 41972 15521 41981 15555
rect 41981 15521 42015 15555
rect 42015 15521 42024 15555
rect 41972 15512 42024 15521
rect 43260 15512 43312 15564
rect 40868 15444 40920 15496
rect 43444 15444 43496 15496
rect 43996 15444 44048 15496
rect 47584 15512 47636 15564
rect 47124 15487 47176 15496
rect 47124 15453 47133 15487
rect 47133 15453 47167 15487
rect 47167 15453 47176 15487
rect 47124 15444 47176 15453
rect 53104 15444 53156 15496
rect 37648 15419 37700 15428
rect 37648 15385 37657 15419
rect 37657 15385 37691 15419
rect 37691 15385 37700 15419
rect 37648 15376 37700 15385
rect 47952 15376 48004 15428
rect 53012 15376 53064 15428
rect 37832 15351 37884 15360
rect 37832 15317 37841 15351
rect 37841 15317 37875 15351
rect 37875 15317 37884 15351
rect 37832 15308 37884 15317
rect 41236 15308 41288 15360
rect 44364 15308 44416 15360
rect 46940 15351 46992 15360
rect 46940 15317 46949 15351
rect 46949 15317 46983 15351
rect 46983 15317 46992 15351
rect 46940 15308 46992 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 1952 15104 2004 15156
rect 4252 15104 4304 15156
rect 4804 15104 4856 15156
rect 5632 15147 5684 15156
rect 5632 15113 5641 15147
rect 5641 15113 5675 15147
rect 5675 15113 5684 15147
rect 5632 15104 5684 15113
rect 8208 15104 8260 15156
rect 9496 15104 9548 15156
rect 12072 15147 12124 15156
rect 12072 15113 12081 15147
rect 12081 15113 12115 15147
rect 12115 15113 12124 15147
rect 12072 15104 12124 15113
rect 12164 15104 12216 15156
rect 2596 15036 2648 15088
rect 2688 14968 2740 15020
rect 3792 14968 3844 15020
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 5080 14968 5132 15020
rect 7564 14968 7616 15020
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 7012 14900 7064 14952
rect 12164 14900 12216 14952
rect 12440 14900 12492 14952
rect 13544 15036 13596 15088
rect 17960 15104 18012 15156
rect 21824 15104 21876 15156
rect 22100 15104 22152 15156
rect 27160 15104 27212 15156
rect 30380 15104 30432 15156
rect 36728 15104 36780 15156
rect 37648 15104 37700 15156
rect 41236 15104 41288 15156
rect 47032 15104 47084 15156
rect 53012 15147 53064 15156
rect 53012 15113 53021 15147
rect 53021 15113 53055 15147
rect 53055 15113 53064 15147
rect 53012 15104 53064 15113
rect 13360 14968 13412 15020
rect 21640 15036 21692 15088
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 8576 14832 8628 14884
rect 10140 14832 10192 14884
rect 16580 14968 16632 15020
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 18696 14968 18748 15020
rect 20904 14968 20956 15020
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 18144 14900 18196 14952
rect 18328 14943 18380 14952
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 18788 14900 18840 14952
rect 21640 14900 21692 14952
rect 30932 15079 30984 15088
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 22468 14968 22520 15020
rect 23296 14968 23348 15020
rect 27068 14968 27120 15020
rect 30932 15045 30941 15079
rect 30941 15045 30975 15079
rect 30975 15045 30984 15079
rect 30932 15036 30984 15045
rect 26608 14900 26660 14952
rect 27436 15011 27488 15020
rect 27436 14977 27450 15011
rect 27450 14977 27484 15011
rect 27484 14977 27488 15011
rect 27436 14968 27488 14977
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 28264 15011 28316 15020
rect 27620 14968 27672 14977
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 30472 14968 30524 15020
rect 32404 15036 32456 15088
rect 34520 15036 34572 15088
rect 37280 15036 37332 15088
rect 40868 15079 40920 15088
rect 30932 14900 30984 14952
rect 35992 14968 36044 15020
rect 40868 15045 40877 15079
rect 40877 15045 40911 15079
rect 40911 15045 40920 15079
rect 40868 15036 40920 15045
rect 43720 15036 43772 15088
rect 46940 15036 46992 15088
rect 37464 14968 37516 15020
rect 38752 14968 38804 15020
rect 43996 14968 44048 15020
rect 44364 15011 44416 15020
rect 44364 14977 44373 15011
rect 44373 14977 44407 15011
rect 44407 14977 44416 15011
rect 44364 14968 44416 14977
rect 46664 14968 46716 15020
rect 47952 14968 48004 15020
rect 53196 15011 53248 15020
rect 53196 14977 53205 15011
rect 53205 14977 53239 15011
rect 53239 14977 53248 15011
rect 53196 14968 53248 14977
rect 31760 14900 31812 14952
rect 37004 14900 37056 14952
rect 3516 14764 3568 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 9956 14764 10008 14816
rect 11152 14764 11204 14816
rect 13268 14764 13320 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 15200 14764 15252 14816
rect 18788 14764 18840 14816
rect 21640 14764 21692 14816
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22284 14832 22336 14884
rect 32312 14832 32364 14884
rect 27896 14764 27948 14816
rect 28080 14807 28132 14816
rect 28080 14773 28089 14807
rect 28089 14773 28123 14807
rect 28123 14773 28132 14807
rect 28080 14764 28132 14773
rect 28172 14764 28224 14816
rect 33324 14764 33376 14816
rect 43260 14807 43312 14816
rect 43260 14773 43269 14807
rect 43269 14773 43303 14807
rect 43303 14773 43312 14807
rect 43260 14764 43312 14773
rect 44180 14764 44232 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2688 14603 2740 14612
rect 2688 14569 2697 14603
rect 2697 14569 2731 14603
rect 2731 14569 2740 14603
rect 2688 14560 2740 14569
rect 5080 14560 5132 14612
rect 9588 14560 9640 14612
rect 10784 14560 10836 14612
rect 13268 14560 13320 14612
rect 15476 14560 15528 14612
rect 16028 14560 16080 14612
rect 16120 14560 16172 14612
rect 16580 14603 16632 14612
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 11612 14492 11664 14544
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 18144 14603 18196 14612
rect 18144 14569 18153 14603
rect 18153 14569 18187 14603
rect 18187 14569 18196 14603
rect 18144 14560 18196 14569
rect 18328 14560 18380 14612
rect 25964 14560 26016 14612
rect 27436 14560 27488 14612
rect 27896 14560 27948 14612
rect 31208 14560 31260 14612
rect 31392 14560 31444 14612
rect 32404 14560 32456 14612
rect 34060 14560 34112 14612
rect 35900 14560 35952 14612
rect 37372 14603 37424 14612
rect 37372 14569 37381 14603
rect 37381 14569 37415 14603
rect 37415 14569 37424 14603
rect 37372 14560 37424 14569
rect 37464 14603 37516 14612
rect 37464 14569 37473 14603
rect 37473 14569 37507 14603
rect 37507 14569 37516 14603
rect 37464 14560 37516 14569
rect 38660 14560 38712 14612
rect 43444 14560 43496 14612
rect 2872 14399 2924 14408
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 6736 14356 6788 14408
rect 7656 14424 7708 14476
rect 14372 14467 14424 14476
rect 5632 14220 5684 14272
rect 7472 14220 7524 14272
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 10508 14399 10560 14408
rect 7748 14356 7800 14365
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 8208 14288 8260 14340
rect 9496 14288 9548 14340
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 15016 14356 15068 14408
rect 15660 14356 15712 14408
rect 9588 14220 9640 14272
rect 10784 14220 10836 14272
rect 16028 14288 16080 14340
rect 18236 14424 18288 14476
rect 23204 14424 23256 14476
rect 25044 14424 25096 14476
rect 26516 14424 26568 14476
rect 28264 14492 28316 14544
rect 31668 14492 31720 14544
rect 18328 14399 18380 14408
rect 18328 14365 18337 14399
rect 18337 14365 18371 14399
rect 18371 14365 18380 14399
rect 18328 14356 18380 14365
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 21364 14356 21416 14408
rect 22928 14356 22980 14408
rect 23020 14356 23072 14408
rect 25872 14356 25924 14408
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 26608 14356 26660 14365
rect 27252 14399 27304 14408
rect 11980 14220 12032 14272
rect 20260 14288 20312 14340
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 22192 14288 22244 14340
rect 27252 14365 27261 14399
rect 27261 14365 27295 14399
rect 27295 14365 27304 14399
rect 27252 14356 27304 14365
rect 30380 14424 30432 14476
rect 31024 14467 31076 14476
rect 31024 14433 31033 14467
rect 31033 14433 31067 14467
rect 31067 14433 31076 14467
rect 31024 14424 31076 14433
rect 39120 14492 39172 14544
rect 43720 14535 43772 14544
rect 43720 14501 43729 14535
rect 43729 14501 43763 14535
rect 43763 14501 43772 14535
rect 43720 14492 43772 14501
rect 34060 14424 34112 14476
rect 34244 14424 34296 14476
rect 28080 14356 28132 14408
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 31116 14356 31168 14408
rect 31392 14356 31444 14408
rect 31668 14356 31720 14408
rect 33600 14356 33652 14408
rect 36360 14356 36412 14408
rect 36728 14356 36780 14408
rect 37004 14399 37056 14408
rect 37004 14365 37013 14399
rect 37013 14365 37047 14399
rect 37047 14365 37056 14399
rect 37004 14356 37056 14365
rect 37924 14424 37976 14476
rect 38476 14424 38528 14476
rect 43260 14424 43312 14476
rect 28724 14288 28776 14340
rect 28816 14288 28868 14340
rect 32772 14288 32824 14340
rect 27068 14220 27120 14272
rect 28264 14220 28316 14272
rect 30380 14220 30432 14272
rect 31024 14220 31076 14272
rect 35808 14288 35860 14340
rect 40868 14356 40920 14408
rect 44456 14356 44508 14408
rect 48412 14356 48464 14408
rect 33876 14220 33928 14272
rect 46296 14288 46348 14340
rect 50620 14288 50672 14340
rect 54024 14356 54076 14408
rect 54576 14288 54628 14340
rect 36176 14220 36228 14272
rect 37832 14220 37884 14272
rect 41052 14220 41104 14272
rect 47952 14263 48004 14272
rect 47952 14229 47961 14263
rect 47961 14229 47995 14263
rect 47995 14229 48004 14263
rect 47952 14220 48004 14229
rect 50160 14220 50212 14272
rect 53748 14263 53800 14272
rect 53748 14229 53757 14263
rect 53757 14229 53791 14263
rect 53791 14229 53800 14263
rect 53748 14220 53800 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 12440 14016 12492 14068
rect 13544 14016 13596 14068
rect 15476 14016 15528 14068
rect 15660 14016 15712 14068
rect 21364 14016 21416 14068
rect 23020 14016 23072 14068
rect 23204 14059 23256 14068
rect 23204 14025 23213 14059
rect 23213 14025 23247 14059
rect 23247 14025 23256 14059
rect 23204 14016 23256 14025
rect 24400 14016 24452 14068
rect 24492 14016 24544 14068
rect 28816 14016 28868 14068
rect 6092 13948 6144 14000
rect 7748 13948 7800 14000
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 5172 13880 5224 13932
rect 7472 13880 7524 13932
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 11520 13948 11572 14000
rect 11612 13948 11664 14000
rect 16304 13948 16356 14000
rect 21456 13948 21508 14000
rect 27988 13991 28040 14000
rect 27988 13957 27997 13991
rect 27997 13957 28031 13991
rect 28031 13957 28040 13991
rect 27988 13948 28040 13957
rect 30380 13948 30432 14000
rect 30656 14016 30708 14068
rect 31392 14016 31444 14068
rect 32772 14016 32824 14068
rect 46664 14059 46716 14068
rect 40316 13948 40368 14000
rect 40408 13948 40460 14000
rect 3056 13812 3108 13864
rect 7012 13812 7064 13864
rect 10508 13880 10560 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 20260 13880 20312 13932
rect 21916 13880 21968 13932
rect 23940 13880 23992 13932
rect 27896 13880 27948 13932
rect 28724 13880 28776 13932
rect 30288 13880 30340 13932
rect 32128 13923 32180 13932
rect 32128 13889 32137 13923
rect 32137 13889 32171 13923
rect 32171 13889 32180 13923
rect 32128 13880 32180 13889
rect 33692 13923 33744 13932
rect 33692 13889 33701 13923
rect 33701 13889 33735 13923
rect 33735 13889 33744 13923
rect 33692 13880 33744 13889
rect 34244 13880 34296 13932
rect 34796 13923 34848 13932
rect 34796 13889 34830 13923
rect 34830 13889 34848 13923
rect 34796 13880 34848 13889
rect 35900 13880 35952 13932
rect 36728 13923 36780 13932
rect 36728 13889 36737 13923
rect 36737 13889 36771 13923
rect 36771 13889 36780 13923
rect 36728 13880 36780 13889
rect 13084 13812 13136 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13452 13812 13504 13864
rect 15844 13812 15896 13864
rect 16212 13812 16264 13864
rect 26332 13812 26384 13864
rect 27252 13812 27304 13864
rect 29276 13812 29328 13864
rect 30196 13855 30248 13864
rect 30196 13821 30205 13855
rect 30205 13821 30239 13855
rect 30239 13821 30248 13855
rect 30196 13812 30248 13821
rect 34520 13855 34572 13864
rect 34520 13821 34529 13855
rect 34529 13821 34563 13855
rect 34563 13821 34572 13855
rect 34520 13812 34572 13821
rect 38752 13812 38804 13864
rect 40040 13812 40092 13864
rect 41052 13923 41104 13932
rect 41052 13889 41061 13923
rect 41061 13889 41095 13923
rect 41095 13889 41104 13923
rect 41052 13880 41104 13889
rect 46664 14025 46673 14059
rect 46673 14025 46707 14059
rect 46707 14025 46716 14059
rect 46664 14016 46716 14025
rect 50620 14059 50672 14068
rect 50620 14025 50629 14059
rect 50629 14025 50663 14059
rect 50663 14025 50672 14059
rect 50620 14016 50672 14025
rect 44456 13948 44508 14000
rect 45008 13880 45060 13932
rect 53196 13948 53248 14000
rect 53748 13948 53800 14000
rect 50528 13923 50580 13932
rect 50528 13889 50537 13923
rect 50537 13889 50571 13923
rect 50571 13889 50580 13923
rect 50528 13880 50580 13889
rect 50620 13880 50672 13932
rect 1860 13744 1912 13796
rect 17224 13744 17276 13796
rect 17316 13744 17368 13796
rect 21640 13744 21692 13796
rect 25872 13744 25924 13796
rect 29000 13744 29052 13796
rect 36544 13744 36596 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 3056 13676 3108 13728
rect 11704 13676 11756 13728
rect 12348 13676 12400 13728
rect 13820 13676 13872 13728
rect 18144 13676 18196 13728
rect 19248 13676 19300 13728
rect 20812 13676 20864 13728
rect 21824 13676 21876 13728
rect 25688 13676 25740 13728
rect 26056 13676 26108 13728
rect 27988 13676 28040 13728
rect 34244 13676 34296 13728
rect 35900 13719 35952 13728
rect 35900 13685 35909 13719
rect 35909 13685 35943 13719
rect 35943 13685 35952 13719
rect 35900 13676 35952 13685
rect 41420 13812 41472 13864
rect 44364 13812 44416 13864
rect 47952 13812 48004 13864
rect 52644 13812 52696 13864
rect 53104 13812 53156 13864
rect 45468 13676 45520 13728
rect 46204 13719 46256 13728
rect 46204 13685 46213 13719
rect 46213 13685 46247 13719
rect 46247 13685 46256 13719
rect 46204 13676 46256 13685
rect 54116 13676 54168 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7380 13472 7432 13524
rect 12624 13472 12676 13524
rect 17224 13472 17276 13524
rect 22836 13472 22888 13524
rect 25688 13472 25740 13524
rect 5172 13447 5224 13456
rect 5172 13413 5181 13447
rect 5181 13413 5215 13447
rect 5215 13413 5224 13447
rect 5172 13404 5224 13413
rect 7932 13404 7984 13456
rect 8576 13404 8628 13456
rect 10508 13404 10560 13456
rect 18512 13404 18564 13456
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 7564 13336 7616 13388
rect 9496 13336 9548 13388
rect 13268 13336 13320 13388
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 7196 13268 7248 13320
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 2228 13243 2280 13252
rect 2228 13209 2237 13243
rect 2237 13209 2271 13243
rect 2271 13209 2280 13243
rect 2228 13200 2280 13209
rect 7104 13200 7156 13252
rect 7564 13200 7616 13252
rect 9404 13132 9456 13184
rect 9588 13268 9640 13320
rect 17224 13268 17276 13320
rect 17960 13200 18012 13252
rect 20168 13336 20220 13388
rect 26792 13404 26844 13456
rect 29920 13472 29972 13524
rect 30104 13472 30156 13524
rect 30840 13472 30892 13524
rect 32864 13472 32916 13524
rect 33416 13515 33468 13524
rect 33416 13481 33425 13515
rect 33425 13481 33459 13515
rect 33459 13481 33468 13515
rect 33416 13472 33468 13481
rect 34796 13472 34848 13524
rect 36360 13515 36412 13524
rect 36360 13481 36369 13515
rect 36369 13481 36403 13515
rect 36403 13481 36412 13515
rect 36360 13472 36412 13481
rect 36728 13472 36780 13524
rect 37004 13472 37056 13524
rect 44088 13515 44140 13524
rect 32128 13404 32180 13456
rect 34244 13404 34296 13456
rect 36820 13404 36872 13456
rect 21732 13336 21784 13388
rect 19432 13268 19484 13320
rect 20076 13268 20128 13320
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 21456 13268 21508 13320
rect 22100 13268 22152 13320
rect 22836 13268 22888 13320
rect 24676 13268 24728 13320
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 26608 13268 26660 13320
rect 27896 13200 27948 13252
rect 28724 13311 28776 13320
rect 28724 13277 28733 13311
rect 28733 13277 28767 13311
rect 28767 13277 28776 13311
rect 28724 13268 28776 13277
rect 29000 13336 29052 13388
rect 34796 13336 34848 13388
rect 29368 13268 29420 13320
rect 30656 13311 30708 13320
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 32128 13311 32180 13320
rect 32128 13277 32137 13311
rect 32137 13277 32171 13311
rect 32171 13277 32180 13311
rect 32128 13268 32180 13277
rect 36084 13268 36136 13320
rect 28172 13200 28224 13252
rect 33140 13243 33192 13252
rect 33140 13209 33149 13243
rect 33149 13209 33183 13243
rect 33183 13209 33192 13243
rect 33140 13200 33192 13209
rect 35900 13200 35952 13252
rect 36268 13268 36320 13320
rect 36912 13268 36964 13320
rect 39764 13268 39816 13320
rect 40684 13268 40736 13320
rect 44088 13481 44097 13515
rect 44097 13481 44131 13515
rect 44131 13481 44140 13515
rect 44088 13472 44140 13481
rect 44456 13515 44508 13524
rect 44456 13481 44465 13515
rect 44465 13481 44499 13515
rect 44499 13481 44508 13515
rect 44456 13472 44508 13481
rect 46296 13472 46348 13524
rect 50528 13472 50580 13524
rect 54576 13515 54628 13524
rect 54576 13481 54585 13515
rect 54585 13481 54619 13515
rect 54619 13481 54628 13515
rect 54576 13472 54628 13481
rect 45468 13404 45520 13456
rect 41144 13379 41196 13388
rect 41144 13345 41153 13379
rect 41153 13345 41187 13379
rect 41187 13345 41196 13379
rect 41144 13336 41196 13345
rect 44180 13379 44232 13388
rect 44180 13345 44189 13379
rect 44189 13345 44223 13379
rect 44223 13345 44232 13379
rect 44180 13336 44232 13345
rect 41420 13311 41472 13320
rect 41420 13277 41454 13311
rect 41454 13277 41472 13311
rect 41420 13268 41472 13277
rect 44364 13268 44416 13320
rect 46204 13311 46256 13320
rect 46204 13277 46213 13311
rect 46213 13277 46247 13311
rect 46247 13277 46256 13311
rect 46204 13268 46256 13277
rect 48044 13404 48096 13456
rect 49148 13311 49200 13320
rect 49148 13277 49157 13311
rect 49157 13277 49191 13311
rect 49191 13277 49200 13311
rect 49148 13268 49200 13277
rect 50160 13268 50212 13320
rect 54944 13336 54996 13388
rect 50988 13268 51040 13320
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 13912 13132 13964 13184
rect 16120 13132 16172 13184
rect 18696 13132 18748 13184
rect 22928 13132 22980 13184
rect 24400 13132 24452 13184
rect 26516 13132 26568 13184
rect 28356 13132 28408 13184
rect 28908 13132 28960 13184
rect 29276 13132 29328 13184
rect 31668 13132 31720 13184
rect 40408 13175 40460 13184
rect 40408 13141 40417 13175
rect 40417 13141 40451 13175
rect 40451 13141 40460 13175
rect 40408 13132 40460 13141
rect 40960 13132 41012 13184
rect 44640 13200 44692 13252
rect 53748 13311 53800 13320
rect 53748 13277 53757 13311
rect 53757 13277 53791 13311
rect 53791 13277 53800 13311
rect 53748 13268 53800 13277
rect 54116 13200 54168 13252
rect 49240 13175 49292 13184
rect 49240 13141 49249 13175
rect 49249 13141 49283 13175
rect 49283 13141 49292 13175
rect 49240 13132 49292 13141
rect 54024 13132 54076 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 7748 12928 7800 12980
rect 9956 12971 10008 12980
rect 5908 12860 5960 12912
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 17960 12971 18012 12980
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7564 12792 7616 12844
rect 3976 12724 4028 12776
rect 7748 12724 7800 12776
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 10876 12792 10928 12844
rect 12532 12860 12584 12912
rect 15292 12903 15344 12912
rect 15292 12869 15301 12903
rect 15301 12869 15335 12903
rect 15335 12869 15344 12903
rect 15292 12860 15344 12869
rect 10140 12724 10192 12776
rect 13084 12792 13136 12844
rect 16120 12860 16172 12912
rect 17960 12937 17969 12971
rect 17969 12937 18003 12971
rect 18003 12937 18012 12971
rect 17960 12928 18012 12937
rect 18512 12928 18564 12980
rect 18696 12928 18748 12980
rect 19432 12860 19484 12912
rect 19984 12903 20036 12912
rect 19984 12869 19993 12903
rect 19993 12869 20027 12903
rect 20027 12869 20036 12903
rect 19984 12860 20036 12869
rect 20812 12903 20864 12912
rect 20812 12869 20821 12903
rect 20821 12869 20855 12903
rect 20855 12869 20864 12903
rect 20812 12860 20864 12869
rect 21456 12928 21508 12980
rect 24860 12928 24912 12980
rect 27988 12860 28040 12912
rect 28356 12903 28408 12912
rect 28356 12869 28365 12903
rect 28365 12869 28399 12903
rect 28399 12869 28408 12903
rect 28356 12860 28408 12869
rect 18144 12835 18196 12844
rect 18144 12801 18172 12835
rect 18172 12801 18196 12835
rect 18144 12792 18196 12801
rect 19156 12792 19208 12844
rect 26056 12792 26108 12844
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 28264 12835 28316 12844
rect 28264 12801 28271 12835
rect 28271 12801 28316 12835
rect 28264 12792 28316 12801
rect 28448 12835 28500 12844
rect 28448 12801 28457 12835
rect 28457 12801 28491 12835
rect 28491 12801 28500 12835
rect 28448 12792 28500 12801
rect 28724 12792 28776 12844
rect 29276 12928 29328 12980
rect 33140 12928 33192 12980
rect 48044 12971 48096 12980
rect 48044 12937 48053 12971
rect 48053 12937 48087 12971
rect 48087 12937 48096 12971
rect 48044 12928 48096 12937
rect 50988 12971 51040 12980
rect 50988 12937 50997 12971
rect 50997 12937 51031 12971
rect 51031 12937 51040 12971
rect 50988 12928 51040 12937
rect 52644 12928 52696 12980
rect 55864 12928 55916 12980
rect 30104 12860 30156 12912
rect 40408 12860 40460 12912
rect 44640 12903 44692 12912
rect 44640 12869 44649 12903
rect 44649 12869 44683 12903
rect 44683 12869 44692 12903
rect 44640 12860 44692 12869
rect 47860 12860 47912 12912
rect 48228 12860 48280 12912
rect 49240 12860 49292 12912
rect 13268 12724 13320 12776
rect 19248 12724 19300 12776
rect 24400 12767 24452 12776
rect 13452 12656 13504 12708
rect 14372 12656 14424 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2872 12588 2924 12640
rect 9680 12588 9732 12640
rect 10968 12588 11020 12640
rect 13636 12588 13688 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 16304 12656 16356 12708
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 29368 12835 29420 12844
rect 29368 12801 29375 12835
rect 29375 12801 29420 12835
rect 29368 12792 29420 12801
rect 38752 12835 38804 12844
rect 38752 12801 38761 12835
rect 38761 12801 38795 12835
rect 38795 12801 38804 12835
rect 38752 12792 38804 12801
rect 39764 12835 39816 12844
rect 39764 12801 39773 12835
rect 39773 12801 39807 12835
rect 39807 12801 39816 12835
rect 39764 12792 39816 12801
rect 40960 12835 41012 12844
rect 40960 12801 40969 12835
rect 40969 12801 41003 12835
rect 41003 12801 41012 12835
rect 40960 12792 41012 12801
rect 44088 12835 44140 12844
rect 40868 12724 40920 12776
rect 44088 12801 44097 12835
rect 44097 12801 44131 12835
rect 44131 12801 44140 12835
rect 44088 12792 44140 12801
rect 44180 12792 44232 12844
rect 45652 12792 45704 12844
rect 50804 12835 50856 12844
rect 50804 12801 50813 12835
rect 50813 12801 50847 12835
rect 50847 12801 50856 12835
rect 50804 12792 50856 12801
rect 53840 12835 53892 12844
rect 17224 12588 17276 12640
rect 24676 12656 24728 12708
rect 28816 12656 28868 12708
rect 39212 12656 39264 12708
rect 48412 12724 48464 12776
rect 44272 12656 44324 12708
rect 45744 12656 45796 12708
rect 46664 12656 46716 12708
rect 50896 12724 50948 12776
rect 53840 12801 53849 12835
rect 53849 12801 53883 12835
rect 53883 12801 53892 12835
rect 53840 12792 53892 12801
rect 54208 12792 54260 12844
rect 55496 12860 55548 12912
rect 55312 12792 55364 12844
rect 54024 12724 54076 12776
rect 54944 12767 54996 12776
rect 54944 12733 54953 12767
rect 54953 12733 54987 12767
rect 54987 12733 54996 12767
rect 54944 12724 54996 12733
rect 55864 12767 55916 12776
rect 55864 12733 55873 12767
rect 55873 12733 55907 12767
rect 55907 12733 55916 12767
rect 55864 12724 55916 12733
rect 21180 12631 21232 12640
rect 21180 12597 21189 12631
rect 21189 12597 21223 12631
rect 21223 12597 21232 12631
rect 21180 12588 21232 12597
rect 22100 12588 22152 12640
rect 22560 12588 22612 12640
rect 26148 12588 26200 12640
rect 27436 12588 27488 12640
rect 28632 12588 28684 12640
rect 28954 12588 29006 12640
rect 31116 12588 31168 12640
rect 37280 12588 37332 12640
rect 39856 12588 39908 12640
rect 45560 12588 45612 12640
rect 53932 12631 53984 12640
rect 53932 12597 53941 12631
rect 53941 12597 53975 12631
rect 53975 12597 53984 12631
rect 53932 12588 53984 12597
rect 54760 12631 54812 12640
rect 54760 12597 54769 12631
rect 54769 12597 54803 12631
rect 54803 12597 54812 12631
rect 54760 12588 54812 12597
rect 55220 12588 55272 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2688 12384 2740 12436
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 21916 12427 21968 12436
rect 4068 12316 4120 12368
rect 7472 12316 7524 12368
rect 2596 12248 2648 12300
rect 1400 12180 1452 12232
rect 4620 12180 4672 12232
rect 5448 12112 5500 12164
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 10232 12316 10284 12368
rect 10784 12316 10836 12368
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 32220 12384 32272 12436
rect 32496 12384 32548 12436
rect 22744 12359 22796 12368
rect 22744 12325 22753 12359
rect 22753 12325 22787 12359
rect 22787 12325 22796 12359
rect 22744 12316 22796 12325
rect 24124 12316 24176 12368
rect 9404 12248 9456 12257
rect 11612 12248 11664 12300
rect 17224 12248 17276 12300
rect 19432 12248 19484 12300
rect 21456 12248 21508 12300
rect 22100 12248 22152 12300
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 7196 12180 7248 12232
rect 7748 12180 7800 12232
rect 7380 12112 7432 12164
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 6736 12044 6788 12096
rect 9036 12180 9088 12232
rect 9220 12180 9272 12232
rect 9496 12180 9548 12232
rect 10508 12180 10560 12232
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 14280 12180 14332 12232
rect 16672 12180 16724 12232
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 18420 12180 18472 12232
rect 21272 12180 21324 12232
rect 22928 12223 22980 12232
rect 22928 12189 22937 12223
rect 22937 12189 22971 12223
rect 22971 12189 22980 12223
rect 22928 12180 22980 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 25320 12180 25372 12232
rect 26148 12180 26200 12232
rect 8852 12044 8904 12096
rect 15108 12112 15160 12164
rect 15936 12112 15988 12164
rect 22652 12112 22704 12164
rect 23572 12112 23624 12164
rect 9404 12044 9456 12096
rect 9680 12044 9732 12096
rect 10416 12044 10468 12096
rect 13544 12044 13596 12096
rect 15292 12044 15344 12096
rect 16396 12044 16448 12096
rect 22100 12044 22152 12096
rect 23020 12044 23072 12096
rect 25596 12044 25648 12096
rect 26424 12223 26476 12232
rect 26424 12189 26438 12223
rect 26438 12189 26472 12223
rect 26472 12189 26476 12223
rect 26424 12180 26476 12189
rect 27252 12112 27304 12164
rect 26516 12044 26568 12096
rect 30196 12248 30248 12300
rect 34520 12384 34572 12436
rect 36084 12384 36136 12436
rect 40316 12384 40368 12436
rect 44272 12384 44324 12436
rect 49148 12384 49200 12436
rect 28172 12180 28224 12232
rect 32128 12180 32180 12232
rect 32312 12223 32364 12232
rect 32312 12189 32321 12223
rect 32321 12189 32355 12223
rect 32355 12189 32364 12223
rect 32312 12180 32364 12189
rect 33968 12180 34020 12232
rect 36544 12180 36596 12232
rect 31760 12155 31812 12164
rect 31760 12121 31769 12155
rect 31769 12121 31803 12155
rect 31803 12121 31812 12155
rect 31760 12112 31812 12121
rect 34704 12112 34756 12164
rect 37096 12180 37148 12232
rect 37280 12180 37332 12232
rect 39856 12223 39908 12232
rect 33692 12044 33744 12096
rect 38476 12112 38528 12164
rect 39856 12189 39871 12223
rect 39871 12189 39905 12223
rect 39905 12189 39908 12223
rect 40684 12223 40736 12232
rect 39856 12180 39908 12189
rect 40684 12189 40693 12223
rect 40693 12189 40727 12223
rect 40727 12189 40736 12223
rect 40684 12180 40736 12189
rect 44180 12316 44232 12368
rect 42432 12248 42484 12300
rect 44916 12180 44968 12232
rect 37372 12044 37424 12096
rect 37464 12087 37516 12096
rect 37464 12053 37473 12087
rect 37473 12053 37507 12087
rect 37507 12053 37516 12087
rect 40868 12112 40920 12164
rect 43260 12155 43312 12164
rect 43260 12121 43269 12155
rect 43269 12121 43303 12155
rect 43303 12121 43312 12155
rect 44272 12155 44324 12164
rect 43260 12112 43312 12121
rect 37464 12044 37516 12053
rect 41144 12044 41196 12096
rect 42432 12044 42484 12096
rect 43720 12087 43772 12096
rect 43720 12053 43729 12087
rect 43729 12053 43763 12087
rect 43763 12053 43772 12087
rect 43720 12044 43772 12053
rect 44272 12121 44281 12155
rect 44281 12121 44315 12155
rect 44315 12121 44324 12155
rect 44272 12112 44324 12121
rect 44364 12087 44416 12096
rect 44364 12053 44373 12087
rect 44373 12053 44407 12087
rect 44407 12053 44416 12087
rect 44364 12044 44416 12053
rect 48596 12248 48648 12300
rect 45560 12223 45612 12232
rect 45560 12189 45594 12223
rect 45594 12189 45612 12223
rect 45560 12180 45612 12189
rect 49700 12180 49752 12232
rect 50620 12427 50672 12436
rect 50620 12393 50629 12427
rect 50629 12393 50663 12427
rect 50663 12393 50672 12427
rect 55312 12427 55364 12436
rect 50620 12384 50672 12393
rect 50896 12316 50948 12368
rect 55312 12393 55321 12427
rect 55321 12393 55355 12427
rect 55355 12393 55364 12427
rect 55312 12384 55364 12393
rect 53748 12316 53800 12368
rect 53840 12316 53892 12368
rect 53748 12223 53800 12232
rect 50160 12112 50212 12164
rect 53748 12189 53757 12223
rect 53757 12189 53791 12223
rect 53791 12189 53800 12223
rect 53748 12180 53800 12189
rect 54024 12223 54076 12232
rect 54024 12189 54033 12223
rect 54033 12189 54067 12223
rect 54067 12189 54076 12223
rect 54024 12180 54076 12189
rect 54208 12180 54260 12232
rect 54760 12180 54812 12232
rect 54116 12112 54168 12164
rect 55220 12112 55272 12164
rect 55496 12155 55548 12164
rect 55496 12121 55505 12155
rect 55505 12121 55539 12155
rect 55539 12121 55548 12155
rect 55496 12112 55548 12121
rect 45560 12044 45612 12096
rect 49700 12044 49752 12096
rect 50804 12044 50856 12096
rect 50988 12044 51040 12096
rect 52000 12087 52052 12096
rect 52000 12053 52009 12087
rect 52009 12053 52043 12087
rect 52043 12053 52052 12087
rect 52000 12044 52052 12053
rect 53564 12087 53616 12096
rect 53564 12053 53573 12087
rect 53573 12053 53607 12087
rect 53607 12053 53616 12087
rect 53564 12044 53616 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2688 11840 2740 11892
rect 7104 11840 7156 11892
rect 8760 11840 8812 11892
rect 13820 11840 13872 11892
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15384 11840 15436 11892
rect 20352 11840 20404 11892
rect 21272 11840 21324 11892
rect 25320 11840 25372 11892
rect 25964 11883 26016 11892
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 2044 11704 2096 11756
rect 3792 11772 3844 11824
rect 6736 11772 6788 11824
rect 7472 11772 7524 11824
rect 7656 11772 7708 11824
rect 2872 11747 2924 11756
rect 2872 11713 2906 11747
rect 2906 11713 2924 11747
rect 2872 11704 2924 11713
rect 6276 11704 6328 11756
rect 7196 11704 7248 11756
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 13544 11772 13596 11824
rect 13728 11815 13780 11824
rect 13728 11781 13737 11815
rect 13737 11781 13771 11815
rect 13771 11781 13780 11815
rect 13728 11772 13780 11781
rect 6920 11636 6972 11688
rect 7840 11636 7892 11688
rect 8760 11704 8812 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 10508 11704 10560 11756
rect 10600 11704 10652 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 11980 11747 12032 11756
rect 11980 11713 11994 11747
rect 11994 11713 12028 11747
rect 12028 11713 12032 11747
rect 11980 11704 12032 11713
rect 12532 11704 12584 11756
rect 12624 11636 12676 11688
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15660 11704 15712 11756
rect 18144 11704 18196 11756
rect 18604 11704 18656 11756
rect 20904 11704 20956 11756
rect 15752 11636 15804 11688
rect 17408 11679 17460 11688
rect 17408 11645 17417 11679
rect 17417 11645 17451 11679
rect 17451 11645 17460 11679
rect 17408 11636 17460 11645
rect 17684 11679 17736 11688
rect 5356 11568 5408 11620
rect 2504 11500 2556 11552
rect 6460 11500 6512 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 10416 11500 10468 11552
rect 17316 11500 17368 11552
rect 17684 11645 17693 11679
rect 17693 11645 17727 11679
rect 17727 11645 17736 11679
rect 17684 11636 17736 11645
rect 17960 11636 18012 11688
rect 18236 11679 18288 11688
rect 18236 11645 18245 11679
rect 18245 11645 18279 11679
rect 18279 11645 18288 11679
rect 18236 11636 18288 11645
rect 21456 11704 21508 11756
rect 21824 11747 21876 11756
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 22744 11772 22796 11824
rect 25228 11772 25280 11824
rect 25596 11815 25648 11824
rect 25596 11781 25605 11815
rect 25605 11781 25639 11815
rect 25639 11781 25648 11815
rect 25596 11772 25648 11781
rect 25964 11849 25973 11883
rect 25973 11849 26007 11883
rect 26007 11849 26016 11883
rect 25964 11840 26016 11849
rect 26056 11840 26108 11892
rect 30472 11840 30524 11892
rect 28080 11772 28132 11824
rect 29920 11815 29972 11824
rect 29920 11781 29929 11815
rect 29929 11781 29963 11815
rect 29963 11781 29972 11815
rect 29920 11772 29972 11781
rect 23020 11704 23072 11756
rect 25320 11747 25372 11756
rect 25320 11713 25329 11747
rect 25329 11713 25363 11747
rect 25363 11713 25372 11747
rect 25320 11704 25372 11713
rect 25688 11747 25740 11756
rect 17592 11568 17644 11620
rect 21640 11636 21692 11688
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 25780 11747 25832 11756
rect 25780 11713 25794 11747
rect 25794 11713 25828 11747
rect 25828 11713 25832 11747
rect 25780 11704 25832 11713
rect 26148 11704 26200 11756
rect 27344 11704 27396 11756
rect 27436 11704 27488 11756
rect 30656 11772 30708 11824
rect 33968 11815 34020 11824
rect 33968 11781 33977 11815
rect 33977 11781 34011 11815
rect 34011 11781 34020 11815
rect 33968 11772 34020 11781
rect 35992 11772 36044 11824
rect 32128 11747 32180 11756
rect 32128 11713 32137 11747
rect 32137 11713 32171 11747
rect 32171 11713 32180 11747
rect 32128 11704 32180 11713
rect 34520 11704 34572 11756
rect 35348 11704 35400 11756
rect 28540 11679 28592 11688
rect 28540 11645 28549 11679
rect 28549 11645 28583 11679
rect 28583 11645 28592 11679
rect 28540 11636 28592 11645
rect 23204 11611 23256 11620
rect 23204 11577 23213 11611
rect 23213 11577 23247 11611
rect 23247 11577 23256 11611
rect 23204 11568 23256 11577
rect 23296 11568 23348 11620
rect 26056 11568 26108 11620
rect 28724 11568 28776 11620
rect 32312 11636 32364 11688
rect 37372 11772 37424 11824
rect 37096 11704 37148 11756
rect 39212 11747 39264 11756
rect 38384 11636 38436 11688
rect 39212 11713 39221 11747
rect 39221 11713 39255 11747
rect 39255 11713 39264 11747
rect 39212 11704 39264 11713
rect 39856 11704 39908 11756
rect 40224 11747 40276 11756
rect 40224 11713 40233 11747
rect 40233 11713 40267 11747
rect 40267 11713 40276 11747
rect 40224 11704 40276 11713
rect 40316 11747 40368 11756
rect 40316 11713 40325 11747
rect 40325 11713 40359 11747
rect 40359 11713 40368 11747
rect 44824 11772 44876 11824
rect 45744 11772 45796 11824
rect 48504 11815 48556 11824
rect 48504 11781 48513 11815
rect 48513 11781 48547 11815
rect 48547 11781 48556 11815
rect 48504 11772 48556 11781
rect 40316 11704 40368 11713
rect 41493 11747 41545 11756
rect 41493 11713 41518 11747
rect 41518 11713 41545 11747
rect 41493 11704 41545 11713
rect 41052 11636 41104 11688
rect 41144 11679 41196 11688
rect 41144 11645 41153 11679
rect 41153 11645 41187 11679
rect 41187 11645 41196 11679
rect 41144 11636 41196 11645
rect 23112 11500 23164 11552
rect 25780 11500 25832 11552
rect 26424 11500 26476 11552
rect 30288 11500 30340 11552
rect 32220 11543 32272 11552
rect 32220 11509 32229 11543
rect 32229 11509 32263 11543
rect 32263 11509 32272 11543
rect 32220 11500 32272 11509
rect 32956 11500 33008 11552
rect 33324 11500 33376 11552
rect 33876 11500 33928 11552
rect 36360 11568 36412 11620
rect 41972 11704 42024 11756
rect 42524 11704 42576 11756
rect 49700 11704 49752 11756
rect 51540 11772 51592 11824
rect 53564 11840 53616 11892
rect 53656 11772 53708 11824
rect 54024 11704 54076 11756
rect 55864 11747 55916 11756
rect 55864 11713 55873 11747
rect 55873 11713 55907 11747
rect 55907 11713 55916 11747
rect 55864 11704 55916 11713
rect 42432 11679 42484 11688
rect 42432 11645 42441 11679
rect 42441 11645 42475 11679
rect 42475 11645 42484 11679
rect 42432 11636 42484 11645
rect 44088 11568 44140 11620
rect 45652 11568 45704 11620
rect 35532 11500 35584 11552
rect 36084 11500 36136 11552
rect 37556 11500 37608 11552
rect 37740 11500 37792 11552
rect 44916 11543 44968 11552
rect 44916 11509 44925 11543
rect 44925 11509 44959 11543
rect 44959 11509 44968 11543
rect 44916 11500 44968 11509
rect 48228 11500 48280 11552
rect 48596 11500 48648 11552
rect 52000 11568 52052 11620
rect 51816 11543 51868 11552
rect 51816 11509 51825 11543
rect 51825 11509 51859 11543
rect 51859 11509 51868 11543
rect 51816 11500 51868 11509
rect 53932 11543 53984 11552
rect 53932 11509 53941 11543
rect 53941 11509 53975 11543
rect 53975 11509 53984 11543
rect 53932 11500 53984 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 10600 11339 10652 11348
rect 10600 11305 10609 11339
rect 10609 11305 10643 11339
rect 10643 11305 10652 11339
rect 10600 11296 10652 11305
rect 11796 11296 11848 11348
rect 15476 11296 15528 11348
rect 17408 11296 17460 11348
rect 1584 11271 1636 11280
rect 1584 11237 1593 11271
rect 1593 11237 1627 11271
rect 1627 11237 1636 11271
rect 1584 11228 1636 11237
rect 6828 11228 6880 11280
rect 7196 11228 7248 11280
rect 9772 11228 9824 11280
rect 11060 11228 11112 11280
rect 11612 11271 11664 11280
rect 11612 11237 11621 11271
rect 11621 11237 11655 11271
rect 11655 11237 11664 11271
rect 11612 11228 11664 11237
rect 4068 11160 4120 11212
rect 7012 11160 7064 11212
rect 7564 11160 7616 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 17316 11228 17368 11280
rect 18052 11160 18104 11212
rect 18328 11203 18380 11212
rect 18328 11169 18337 11203
rect 18337 11169 18371 11203
rect 18371 11169 18380 11203
rect 18328 11160 18380 11169
rect 18604 11160 18656 11212
rect 20904 11296 20956 11348
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22560 11339 22612 11348
rect 22376 11296 22428 11305
rect 22560 11305 22569 11339
rect 22569 11305 22603 11339
rect 22603 11305 22612 11339
rect 22560 11296 22612 11305
rect 23112 11296 23164 11348
rect 25228 11296 25280 11348
rect 30656 11296 30708 11348
rect 32312 11296 32364 11348
rect 33600 11296 33652 11348
rect 35348 11296 35400 11348
rect 35532 11339 35584 11348
rect 35532 11305 35541 11339
rect 35541 11305 35575 11339
rect 35575 11305 35584 11339
rect 35532 11296 35584 11305
rect 35716 11296 35768 11348
rect 38752 11296 38804 11348
rect 40224 11296 40276 11348
rect 47676 11296 47728 11348
rect 20352 11228 20404 11280
rect 22192 11228 22244 11280
rect 22284 11228 22336 11280
rect 23204 11228 23256 11280
rect 25504 11228 25556 11280
rect 26148 11228 26200 11280
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 6184 11092 6236 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 6920 11092 6972 11144
rect 7196 11092 7248 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 2320 10956 2372 11008
rect 9956 11024 10008 11076
rect 10048 11024 10100 11076
rect 12072 11092 12124 11144
rect 12348 11092 12400 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15752 11092 15804 11144
rect 18420 11135 18472 11144
rect 10784 10956 10836 11008
rect 11152 10956 11204 11008
rect 13728 11024 13780 11076
rect 14372 11024 14424 11076
rect 16028 11067 16080 11076
rect 16028 11033 16037 11067
rect 16037 11033 16071 11067
rect 16071 11033 16080 11067
rect 16028 11024 16080 11033
rect 16120 11024 16172 11076
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 15016 10999 15068 11008
rect 15016 10965 15025 10999
rect 15025 10965 15059 10999
rect 15059 10965 15068 10999
rect 15016 10956 15068 10965
rect 19524 11067 19576 11076
rect 19524 11033 19558 11067
rect 19558 11033 19576 11067
rect 19524 11024 19576 11033
rect 21548 11024 21600 11076
rect 20628 10999 20680 11008
rect 20628 10965 20637 10999
rect 20637 10965 20671 10999
rect 20671 10965 20680 10999
rect 20628 10956 20680 10965
rect 22284 11024 22336 11076
rect 23020 11092 23072 11144
rect 23388 11135 23440 11144
rect 23388 11101 23395 11135
rect 23395 11101 23440 11135
rect 23388 11092 23440 11101
rect 24492 11135 24544 11144
rect 24492 11101 24501 11135
rect 24501 11101 24535 11135
rect 24535 11101 24544 11135
rect 24492 11092 24544 11101
rect 26332 11135 26384 11144
rect 26332 11101 26341 11135
rect 26341 11101 26375 11135
rect 26375 11101 26384 11135
rect 26332 11092 26384 11101
rect 30196 11160 30248 11212
rect 32956 11135 33008 11144
rect 32956 11101 32965 11135
rect 32965 11101 32999 11135
rect 32999 11101 33008 11135
rect 32956 11092 33008 11101
rect 33324 11092 33376 11144
rect 23296 10956 23348 11008
rect 25780 11024 25832 11076
rect 32128 11024 32180 11076
rect 43260 11228 43312 11280
rect 37556 11160 37608 11212
rect 40868 11160 40920 11212
rect 48596 11296 48648 11348
rect 50896 11339 50948 11348
rect 50896 11305 50905 11339
rect 50905 11305 50939 11339
rect 50939 11305 50948 11339
rect 50896 11296 50948 11305
rect 51540 11296 51592 11348
rect 35716 11092 35768 11144
rect 36268 11135 36320 11144
rect 36268 11101 36277 11135
rect 36277 11101 36311 11135
rect 36311 11101 36320 11135
rect 36268 11092 36320 11101
rect 36360 11135 36412 11144
rect 36360 11101 36369 11135
rect 36369 11101 36403 11135
rect 36403 11101 36412 11135
rect 36544 11135 36596 11144
rect 36360 11092 36412 11101
rect 36544 11101 36553 11135
rect 36553 11101 36587 11135
rect 36587 11101 36596 11135
rect 36544 11092 36596 11101
rect 38476 11092 38528 11144
rect 41512 11092 41564 11144
rect 43720 11092 43772 11144
rect 23664 10956 23716 11008
rect 28448 10956 28500 11008
rect 28908 10956 28960 11008
rect 33048 10999 33100 11008
rect 33048 10965 33057 10999
rect 33057 10965 33091 10999
rect 33091 10965 33100 10999
rect 33048 10956 33100 10965
rect 33232 10956 33284 11008
rect 36084 10999 36136 11008
rect 36084 10965 36093 10999
rect 36093 10965 36127 10999
rect 36127 10965 36136 10999
rect 36084 10956 36136 10965
rect 36360 10956 36412 11008
rect 42432 11024 42484 11076
rect 45560 11024 45612 11076
rect 48320 11024 48372 11076
rect 42984 10956 43036 11008
rect 54392 11092 54444 11144
rect 49884 10956 49936 11008
rect 53104 10956 53156 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 7012 10752 7064 10804
rect 11060 10752 11112 10804
rect 3516 10684 3568 10736
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2320 10659 2372 10668
rect 2320 10625 2354 10659
rect 2354 10625 2372 10659
rect 2320 10616 2372 10625
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 6920 10548 6972 10600
rect 3608 10480 3660 10532
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 7840 10616 7892 10668
rect 7748 10548 7800 10600
rect 10508 10684 10560 10736
rect 10968 10684 11020 10736
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 11704 10616 11756 10668
rect 14096 10684 14148 10736
rect 14372 10684 14424 10736
rect 15016 10684 15068 10736
rect 15200 10684 15252 10736
rect 16396 10684 16448 10736
rect 17684 10684 17736 10736
rect 19432 10684 19484 10736
rect 19524 10727 19576 10736
rect 19524 10693 19533 10727
rect 19533 10693 19567 10727
rect 19567 10693 19576 10727
rect 19524 10684 19576 10693
rect 20628 10684 20680 10736
rect 22376 10752 22428 10804
rect 23388 10752 23440 10804
rect 27344 10752 27396 10804
rect 33048 10752 33100 10804
rect 38752 10752 38804 10804
rect 41972 10752 42024 10804
rect 44548 10752 44600 10804
rect 48504 10752 48556 10804
rect 50804 10752 50856 10804
rect 54392 10795 54444 10804
rect 54392 10761 54401 10795
rect 54401 10761 54435 10795
rect 54435 10761 54444 10795
rect 54392 10752 54444 10761
rect 35532 10684 35584 10736
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 16580 10616 16632 10668
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 14004 10548 14056 10600
rect 19524 10548 19576 10600
rect 7932 10480 7984 10532
rect 10508 10480 10560 10532
rect 10876 10480 10928 10532
rect 16396 10480 16448 10532
rect 19156 10480 19208 10532
rect 27620 10616 27672 10668
rect 32128 10616 32180 10668
rect 36084 10659 36136 10668
rect 36084 10625 36093 10659
rect 36093 10625 36127 10659
rect 36127 10625 36136 10659
rect 36084 10616 36136 10625
rect 36360 10659 36412 10668
rect 36360 10625 36369 10659
rect 36369 10625 36403 10659
rect 36403 10625 36412 10659
rect 36360 10616 36412 10625
rect 48596 10684 48648 10736
rect 49884 10727 49936 10736
rect 30196 10548 30248 10600
rect 42340 10616 42392 10668
rect 49884 10693 49893 10727
rect 49893 10693 49927 10727
rect 49927 10693 49936 10727
rect 49884 10684 49936 10693
rect 49976 10684 50028 10736
rect 53288 10659 53340 10668
rect 53288 10625 53322 10659
rect 53322 10625 53340 10659
rect 53288 10616 53340 10625
rect 48228 10548 48280 10600
rect 3424 10412 3476 10421
rect 7564 10412 7616 10464
rect 7748 10412 7800 10464
rect 11612 10412 11664 10464
rect 16028 10412 16080 10464
rect 31576 10480 31628 10532
rect 33416 10480 33468 10532
rect 52644 10548 52696 10600
rect 32220 10412 32272 10464
rect 35900 10455 35952 10464
rect 35900 10421 35909 10455
rect 35909 10421 35943 10455
rect 35943 10421 35952 10455
rect 35900 10412 35952 10421
rect 43076 10412 43128 10464
rect 50068 10455 50120 10464
rect 50068 10421 50077 10455
rect 50077 10421 50111 10455
rect 50111 10421 50120 10455
rect 50068 10412 50120 10421
rect 50988 10412 51040 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2412 10208 2464 10260
rect 6092 10208 6144 10260
rect 11704 10208 11756 10260
rect 11980 10208 12032 10260
rect 2596 10140 2648 10192
rect 10140 10140 10192 10192
rect 14280 10208 14332 10260
rect 14648 10208 14700 10260
rect 3792 10072 3844 10124
rect 7840 10072 7892 10124
rect 3424 10004 3476 10056
rect 4896 10004 4948 10056
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 16580 10072 16632 10124
rect 7196 10004 7248 10013
rect 11612 10047 11664 10056
rect 11612 10013 11619 10047
rect 11619 10013 11664 10047
rect 11612 10004 11664 10013
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11888 10047 11940 10056
rect 11888 10013 11902 10047
rect 11902 10013 11936 10047
rect 11936 10013 11940 10047
rect 11888 10004 11940 10013
rect 6368 9936 6420 9988
rect 14832 9979 14884 9988
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 6460 9868 6512 9920
rect 10876 9868 10928 9920
rect 14832 9945 14841 9979
rect 14841 9945 14875 9979
rect 14875 9945 14884 9979
rect 14832 9936 14884 9945
rect 15200 9936 15252 9988
rect 18052 10208 18104 10260
rect 34796 10208 34848 10260
rect 36084 10251 36136 10260
rect 36084 10217 36093 10251
rect 36093 10217 36127 10251
rect 36127 10217 36136 10251
rect 36084 10208 36136 10217
rect 36728 10208 36780 10260
rect 42340 10251 42392 10260
rect 42340 10217 42349 10251
rect 42349 10217 42383 10251
rect 42383 10217 42392 10251
rect 42340 10208 42392 10217
rect 47676 10251 47728 10260
rect 47676 10217 47685 10251
rect 47685 10217 47719 10251
rect 47719 10217 47728 10251
rect 47676 10208 47728 10217
rect 49608 10208 49660 10260
rect 53288 10251 53340 10260
rect 53288 10217 53297 10251
rect 53297 10217 53331 10251
rect 53331 10217 53340 10251
rect 53288 10208 53340 10217
rect 26884 10140 26936 10192
rect 31944 10072 31996 10124
rect 18236 10004 18288 10056
rect 19524 10004 19576 10056
rect 21180 10004 21232 10056
rect 26332 10047 26384 10056
rect 26332 10013 26341 10047
rect 26341 10013 26375 10047
rect 26375 10013 26384 10047
rect 26332 10004 26384 10013
rect 36544 10072 36596 10124
rect 32036 9936 32088 9988
rect 17224 9868 17276 9920
rect 18420 9868 18472 9920
rect 25872 9911 25924 9920
rect 25872 9877 25881 9911
rect 25881 9877 25915 9911
rect 25915 9877 25924 9911
rect 25872 9868 25924 9877
rect 27068 9868 27120 9920
rect 31576 9868 31628 9920
rect 33508 10004 33560 10056
rect 34704 10047 34756 10056
rect 34704 10013 34713 10047
rect 34713 10013 34747 10047
rect 34747 10013 34756 10047
rect 34704 10004 34756 10013
rect 37464 10004 37516 10056
rect 39212 10004 39264 10056
rect 40960 10047 41012 10056
rect 40960 10013 40969 10047
rect 40969 10013 41003 10047
rect 41003 10013 41012 10047
rect 40960 10004 41012 10013
rect 42984 10115 43036 10124
rect 42984 10081 42993 10115
rect 42993 10081 43027 10115
rect 43027 10081 43036 10115
rect 42984 10072 43036 10081
rect 45560 10072 45612 10124
rect 52920 10072 52972 10124
rect 41328 10047 41380 10056
rect 41328 10013 41337 10047
rect 41337 10013 41371 10047
rect 41371 10013 41380 10047
rect 41972 10047 42024 10056
rect 41328 10004 41380 10013
rect 41972 10013 41981 10047
rect 41981 10013 42015 10047
rect 42015 10013 42024 10047
rect 41972 10004 42024 10013
rect 42156 10047 42208 10056
rect 42156 10013 42165 10047
rect 42165 10013 42199 10047
rect 42199 10013 42208 10047
rect 42156 10004 42208 10013
rect 43076 10004 43128 10056
rect 32312 9979 32364 9988
rect 32312 9945 32321 9979
rect 32321 9945 32355 9979
rect 32355 9945 32364 9979
rect 32312 9936 32364 9945
rect 33140 9936 33192 9988
rect 36176 9936 36228 9988
rect 32680 9911 32732 9920
rect 32680 9877 32689 9911
rect 32689 9877 32723 9911
rect 32723 9877 32732 9911
rect 32680 9868 32732 9877
rect 35256 9868 35308 9920
rect 35624 9868 35676 9920
rect 36268 9911 36320 9920
rect 36268 9877 36277 9911
rect 36277 9877 36311 9911
rect 36311 9877 36320 9911
rect 36268 9868 36320 9877
rect 38016 9868 38068 9920
rect 45560 9936 45612 9988
rect 53104 10047 53156 10056
rect 53104 10013 53113 10047
rect 53113 10013 53147 10047
rect 53147 10013 53156 10047
rect 53104 10004 53156 10013
rect 53196 10047 53248 10056
rect 53196 10013 53205 10047
rect 53205 10013 53239 10047
rect 53239 10013 53248 10047
rect 53196 10004 53248 10013
rect 53932 9936 53984 9988
rect 41420 9868 41472 9920
rect 41512 9911 41564 9920
rect 41512 9877 41521 9911
rect 41521 9877 41555 9911
rect 41555 9877 41564 9911
rect 41512 9868 41564 9877
rect 43904 9868 43956 9920
rect 47032 9911 47084 9920
rect 47032 9877 47041 9911
rect 47041 9877 47075 9911
rect 47075 9877 47084 9911
rect 47032 9868 47084 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6092 9664 6144 9716
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 11888 9664 11940 9716
rect 3240 9528 3292 9580
rect 7472 9528 7524 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 10600 9596 10652 9648
rect 10968 9596 11020 9648
rect 12348 9664 12400 9716
rect 14832 9664 14884 9716
rect 18236 9664 18288 9716
rect 32036 9664 32088 9716
rect 38660 9664 38712 9716
rect 39212 9664 39264 9716
rect 14556 9596 14608 9648
rect 17132 9596 17184 9648
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 9956 9528 10008 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 14280 9571 14332 9580
rect 13360 9528 13412 9537
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 11704 9460 11756 9512
rect 12992 9460 13044 9512
rect 13912 9460 13964 9512
rect 14648 9460 14700 9512
rect 17040 9460 17092 9512
rect 10600 9392 10652 9444
rect 18236 9571 18288 9580
rect 18236 9537 18245 9571
rect 18245 9537 18279 9571
rect 18279 9537 18288 9571
rect 18236 9528 18288 9537
rect 19340 9528 19392 9580
rect 20076 9528 20128 9580
rect 22376 9571 22428 9580
rect 22376 9537 22410 9571
rect 22410 9537 22428 9571
rect 25872 9596 25924 9648
rect 32404 9596 32456 9648
rect 42156 9664 42208 9716
rect 50712 9707 50764 9716
rect 50712 9673 50721 9707
rect 50721 9673 50755 9707
rect 50755 9673 50764 9707
rect 50712 9664 50764 9673
rect 52644 9664 52696 9716
rect 53564 9664 53616 9716
rect 22376 9528 22428 9537
rect 26884 9528 26936 9580
rect 29552 9528 29604 9580
rect 32680 9528 32732 9580
rect 33140 9571 33192 9580
rect 33140 9537 33149 9571
rect 33149 9537 33183 9571
rect 33183 9537 33192 9571
rect 33140 9528 33192 9537
rect 18052 9460 18104 9512
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 7472 9324 7524 9376
rect 8392 9324 8444 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 9956 9324 10008 9376
rect 10508 9324 10560 9376
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 14372 9324 14424 9376
rect 16856 9324 16908 9376
rect 16948 9324 17000 9376
rect 17684 9392 17736 9444
rect 17776 9324 17828 9376
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 22008 9460 22060 9512
rect 23480 9460 23532 9512
rect 26792 9460 26844 9512
rect 28172 9503 28224 9512
rect 28172 9469 28181 9503
rect 28181 9469 28215 9503
rect 28215 9469 28224 9503
rect 28172 9460 28224 9469
rect 31760 9460 31812 9512
rect 26240 9392 26292 9444
rect 27344 9392 27396 9444
rect 33048 9392 33100 9444
rect 41236 9639 41288 9648
rect 20628 9367 20680 9376
rect 20628 9333 20637 9367
rect 20637 9333 20671 9367
rect 20671 9333 20680 9367
rect 20628 9324 20680 9333
rect 23112 9324 23164 9376
rect 29552 9367 29604 9376
rect 29552 9333 29561 9367
rect 29561 9333 29595 9367
rect 29595 9333 29604 9367
rect 29552 9324 29604 9333
rect 30196 9367 30248 9376
rect 30196 9333 30205 9367
rect 30205 9333 30239 9367
rect 30239 9333 30248 9367
rect 30196 9324 30248 9333
rect 31116 9324 31168 9376
rect 33508 9571 33560 9580
rect 33508 9537 33517 9571
rect 33517 9537 33551 9571
rect 33551 9537 33560 9571
rect 33508 9528 33560 9537
rect 33692 9528 33744 9580
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 36268 9528 36320 9580
rect 37832 9528 37884 9580
rect 41236 9605 41245 9639
rect 41245 9605 41279 9639
rect 41279 9605 41288 9639
rect 41236 9596 41288 9605
rect 45468 9639 45520 9648
rect 45468 9605 45477 9639
rect 45477 9605 45511 9639
rect 45511 9605 45520 9639
rect 45468 9596 45520 9605
rect 33784 9460 33836 9512
rect 38108 9460 38160 9512
rect 40960 9571 41012 9580
rect 40960 9537 40969 9571
rect 40969 9537 41003 9571
rect 41003 9537 41012 9571
rect 40960 9528 41012 9537
rect 41144 9571 41196 9580
rect 41144 9537 41153 9571
rect 41153 9537 41187 9571
rect 41187 9537 41196 9571
rect 41144 9528 41196 9537
rect 41328 9571 41380 9580
rect 41328 9537 41337 9571
rect 41337 9537 41371 9571
rect 41371 9537 41380 9571
rect 41328 9528 41380 9537
rect 41512 9528 41564 9580
rect 33692 9435 33744 9444
rect 33692 9401 33701 9435
rect 33701 9401 33735 9435
rect 33735 9401 33744 9435
rect 33692 9392 33744 9401
rect 35256 9392 35308 9444
rect 35532 9392 35584 9444
rect 38200 9392 38252 9444
rect 34152 9324 34204 9376
rect 35348 9324 35400 9376
rect 36176 9324 36228 9376
rect 37556 9324 37608 9376
rect 38936 9503 38988 9512
rect 38936 9469 38945 9503
rect 38945 9469 38979 9503
rect 38979 9469 38988 9503
rect 38936 9460 38988 9469
rect 41972 9460 42024 9512
rect 47032 9528 47084 9580
rect 48228 9528 48280 9580
rect 49976 9528 50028 9580
rect 51816 9528 51868 9580
rect 53196 9596 53248 9648
rect 39212 9392 39264 9444
rect 48596 9460 48648 9512
rect 49516 9503 49568 9512
rect 49516 9469 49525 9503
rect 49525 9469 49559 9503
rect 49559 9469 49568 9503
rect 49516 9460 49568 9469
rect 49608 9460 49660 9512
rect 45560 9392 45612 9444
rect 50988 9460 51040 9512
rect 54024 9528 54076 9580
rect 53564 9392 53616 9444
rect 41328 9324 41380 9376
rect 45192 9324 45244 9376
rect 53012 9324 53064 9376
rect 53748 9367 53800 9376
rect 53748 9333 53757 9367
rect 53757 9333 53791 9367
rect 53791 9333 53800 9367
rect 53748 9324 53800 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 9496 9120 9548 9172
rect 10968 9163 11020 9172
rect 4344 9052 4396 9104
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11704 9120 11756 9172
rect 17868 9120 17920 9172
rect 20076 9163 20128 9172
rect 16672 9052 16724 9104
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 9496 8984 9548 9036
rect 13912 8984 13964 9036
rect 14648 8984 14700 9036
rect 16580 8984 16632 9036
rect 17316 9052 17368 9104
rect 17132 8984 17184 9036
rect 17776 9027 17828 9036
rect 17776 8993 17785 9027
rect 17785 8993 17819 9027
rect 17819 8993 17828 9027
rect 17776 8984 17828 8993
rect 20076 9129 20085 9163
rect 20085 9129 20119 9163
rect 20119 9129 20128 9163
rect 20076 9120 20128 9129
rect 22376 9120 22428 9172
rect 26332 9120 26384 9172
rect 21364 9052 21416 9104
rect 20628 9027 20680 9036
rect 20628 8993 20637 9027
rect 20637 8993 20671 9027
rect 20671 8993 20680 9027
rect 20628 8984 20680 8993
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 9588 8959 9640 8968
rect 9588 8925 9597 8959
rect 9597 8925 9631 8959
rect 9631 8925 9640 8959
rect 9588 8916 9640 8925
rect 9680 8916 9732 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 14372 8959 14424 8968
rect 11704 8848 11756 8900
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4068 8780 4120 8832
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 10508 8780 10560 8832
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 16764 8959 16816 8968
rect 14556 8916 14608 8925
rect 16764 8925 16773 8959
rect 16773 8925 16807 8959
rect 16807 8925 16816 8959
rect 16764 8916 16816 8925
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 17224 8916 17276 8968
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 23572 9052 23624 9104
rect 23756 9027 23808 9036
rect 21364 8959 21416 8968
rect 14188 8780 14240 8832
rect 15752 8780 15804 8832
rect 20628 8848 20680 8900
rect 20720 8891 20772 8900
rect 20720 8857 20729 8891
rect 20729 8857 20763 8891
rect 20763 8857 20772 8891
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 26056 8984 26108 9036
rect 26884 8984 26936 9036
rect 32312 9120 32364 9172
rect 33508 9120 33560 9172
rect 37556 9120 37608 9172
rect 34336 9052 34388 9104
rect 40040 9120 40092 9172
rect 41420 9120 41472 9172
rect 50712 9120 50764 9172
rect 53012 9120 53064 9172
rect 54024 9163 54076 9172
rect 54024 9129 54033 9163
rect 54033 9129 54067 9163
rect 54067 9129 54076 9163
rect 54024 9120 54076 9129
rect 39120 9052 39172 9104
rect 20720 8848 20772 8857
rect 21732 8848 21784 8900
rect 24584 8916 24636 8968
rect 26240 8916 26292 8968
rect 28172 8916 28224 8968
rect 30012 8959 30064 8968
rect 30012 8925 30021 8959
rect 30021 8925 30055 8959
rect 30055 8925 30064 8959
rect 30012 8916 30064 8925
rect 32404 8984 32456 9036
rect 33692 8984 33744 9036
rect 35900 8984 35952 9036
rect 36820 8984 36872 9036
rect 42156 9052 42208 9104
rect 46940 9052 46992 9104
rect 50160 9095 50212 9104
rect 50160 9061 50169 9095
rect 50169 9061 50203 9095
rect 50203 9061 50212 9095
rect 50160 9052 50212 9061
rect 42524 8984 42576 9036
rect 23112 8891 23164 8900
rect 23112 8857 23121 8891
rect 23121 8857 23155 8891
rect 23155 8857 23164 8891
rect 23112 8848 23164 8857
rect 23204 8891 23256 8900
rect 23204 8857 23213 8891
rect 23213 8857 23247 8891
rect 23247 8857 23256 8891
rect 23204 8848 23256 8857
rect 30932 8848 30984 8900
rect 30840 8780 30892 8832
rect 32496 8848 32548 8900
rect 33600 8848 33652 8900
rect 32036 8780 32088 8832
rect 33968 8823 34020 8832
rect 33968 8789 33977 8823
rect 33977 8789 34011 8823
rect 34011 8789 34020 8823
rect 33968 8780 34020 8789
rect 34152 8959 34204 8968
rect 34152 8925 34161 8959
rect 34161 8925 34195 8959
rect 34195 8925 34204 8959
rect 35348 8959 35400 8968
rect 34152 8916 34204 8925
rect 35348 8925 35357 8959
rect 35357 8925 35391 8959
rect 35391 8925 35400 8959
rect 35348 8916 35400 8925
rect 37924 8959 37976 8968
rect 34336 8848 34388 8900
rect 37924 8925 37933 8959
rect 37933 8925 37967 8959
rect 37967 8925 37976 8959
rect 37924 8916 37976 8925
rect 38016 8916 38068 8968
rect 47032 8984 47084 9036
rect 45192 8959 45244 8968
rect 45192 8925 45201 8959
rect 45201 8925 45235 8959
rect 45235 8925 45244 8959
rect 45192 8916 45244 8925
rect 50068 8916 50120 8968
rect 50712 8916 50764 8968
rect 50988 8916 51040 8968
rect 53288 8916 53340 8968
rect 34704 8780 34756 8832
rect 36544 8780 36596 8832
rect 53656 8891 53708 8900
rect 39304 8823 39356 8832
rect 39304 8789 39313 8823
rect 39313 8789 39347 8823
rect 39347 8789 39356 8823
rect 39304 8780 39356 8789
rect 39396 8780 39448 8832
rect 42156 8823 42208 8832
rect 42156 8789 42165 8823
rect 42165 8789 42199 8823
rect 42199 8789 42208 8823
rect 42156 8780 42208 8789
rect 42616 8780 42668 8832
rect 45008 8823 45060 8832
rect 45008 8789 45017 8823
rect 45017 8789 45051 8823
rect 45051 8789 45060 8823
rect 45008 8780 45060 8789
rect 53656 8857 53665 8891
rect 53665 8857 53699 8891
rect 53699 8857 53708 8891
rect 53656 8848 53708 8857
rect 53748 8848 53800 8900
rect 52920 8780 52972 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 4344 8576 4396 8628
rect 1768 8551 1820 8560
rect 1768 8517 1777 8551
rect 1777 8517 1811 8551
rect 1811 8517 1820 8551
rect 1768 8508 1820 8517
rect 3792 8508 3844 8560
rect 3976 8508 4028 8560
rect 7380 8576 7432 8628
rect 9864 8576 9916 8628
rect 10508 8576 10560 8628
rect 11704 8576 11756 8628
rect 16856 8576 16908 8628
rect 7012 8508 7064 8560
rect 2228 8440 2280 8492
rect 2044 8372 2096 8424
rect 4068 8304 4120 8356
rect 4252 8440 4304 8492
rect 4620 8440 4672 8492
rect 7472 8440 7524 8492
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 13452 8508 13504 8560
rect 14556 8508 14608 8560
rect 9496 8440 9548 8492
rect 8300 8372 8352 8424
rect 10692 8372 10744 8424
rect 12716 8440 12768 8492
rect 13360 8440 13412 8492
rect 13820 8440 13872 8492
rect 14188 8440 14240 8492
rect 14740 8440 14792 8492
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 12992 8304 13044 8313
rect 13084 8304 13136 8356
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 15476 8372 15528 8424
rect 15660 8508 15712 8560
rect 16764 8508 16816 8560
rect 17132 8508 17184 8560
rect 20720 8576 20772 8628
rect 22100 8576 22152 8628
rect 23204 8576 23256 8628
rect 30932 8619 30984 8628
rect 30932 8585 30941 8619
rect 30941 8585 30975 8619
rect 30975 8585 30984 8619
rect 30932 8576 30984 8585
rect 31024 8576 31076 8628
rect 24584 8508 24636 8560
rect 27804 8508 27856 8560
rect 28172 8508 28224 8560
rect 34336 8576 34388 8628
rect 36544 8576 36596 8628
rect 38108 8576 38160 8628
rect 39396 8576 39448 8628
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16212 8440 16264 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 23572 8483 23624 8492
rect 16948 8440 17000 8449
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 23756 8440 23808 8492
rect 16672 8372 16724 8424
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 17040 8415 17092 8424
rect 17040 8381 17049 8415
rect 17049 8381 17083 8415
rect 17083 8381 17092 8415
rect 17040 8372 17092 8381
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17592 8372 17644 8424
rect 23848 8415 23900 8424
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 27528 8440 27580 8492
rect 31116 8483 31168 8492
rect 28080 8372 28132 8424
rect 13452 8236 13504 8288
rect 21364 8304 21416 8356
rect 21732 8304 21784 8356
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 33784 8440 33836 8492
rect 33968 8508 34020 8560
rect 35808 8508 35860 8560
rect 40868 8576 40920 8628
rect 41144 8576 41196 8628
rect 50068 8576 50120 8628
rect 50620 8576 50672 8628
rect 40040 8508 40092 8560
rect 40776 8508 40828 8560
rect 42524 8508 42576 8560
rect 30012 8372 30064 8424
rect 30288 8304 30340 8356
rect 36176 8440 36228 8492
rect 36268 8440 36320 8492
rect 35808 8372 35860 8424
rect 39304 8440 39356 8492
rect 40132 8483 40184 8492
rect 40132 8449 40141 8483
rect 40141 8449 40175 8483
rect 40175 8449 40184 8483
rect 40132 8440 40184 8449
rect 40224 8483 40276 8492
rect 40224 8449 40233 8483
rect 40233 8449 40267 8483
rect 40267 8449 40276 8483
rect 40224 8440 40276 8449
rect 40500 8440 40552 8492
rect 42800 8483 42852 8492
rect 42800 8449 42809 8483
rect 42809 8449 42843 8483
rect 42843 8449 42852 8483
rect 42800 8440 42852 8449
rect 39120 8415 39172 8424
rect 39120 8381 39129 8415
rect 39129 8381 39163 8415
rect 39163 8381 39172 8415
rect 39120 8372 39172 8381
rect 23756 8279 23808 8288
rect 23756 8245 23765 8279
rect 23765 8245 23799 8279
rect 23799 8245 23808 8279
rect 23756 8236 23808 8245
rect 27160 8236 27212 8288
rect 30196 8236 30248 8288
rect 31392 8236 31444 8288
rect 33416 8236 33468 8288
rect 40040 8304 40092 8356
rect 40132 8304 40184 8356
rect 42248 8372 42300 8424
rect 45008 8508 45060 8560
rect 43720 8440 43772 8492
rect 45560 8440 45612 8492
rect 52644 8508 52696 8560
rect 50160 8440 50212 8492
rect 53288 8440 53340 8492
rect 53012 8415 53064 8424
rect 40868 8304 40920 8356
rect 41420 8304 41472 8356
rect 53012 8381 53021 8415
rect 53021 8381 53055 8415
rect 53055 8381 53064 8415
rect 53012 8372 53064 8381
rect 43812 8304 43864 8356
rect 46940 8304 46992 8356
rect 47768 8304 47820 8356
rect 34152 8236 34204 8288
rect 34244 8236 34296 8288
rect 36176 8236 36228 8288
rect 36360 8236 36412 8288
rect 53012 8236 53064 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 16856 8032 16908 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 1952 7828 2004 7880
rect 4620 7828 4672 7880
rect 13728 7964 13780 8016
rect 13084 7896 13136 7948
rect 14556 7896 14608 7948
rect 15936 7896 15988 7948
rect 7472 7828 7524 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10600 7828 10652 7880
rect 11428 7828 11480 7880
rect 13176 7871 13228 7880
rect 9956 7760 10008 7812
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 14188 7828 14240 7880
rect 17224 7964 17276 8016
rect 28080 8032 28132 8084
rect 28724 8032 28776 8084
rect 33048 8075 33100 8084
rect 17684 7939 17736 7948
rect 17684 7905 17693 7939
rect 17693 7905 17727 7939
rect 17727 7905 17736 7939
rect 17684 7896 17736 7905
rect 18420 7896 18472 7948
rect 30288 7964 30340 8016
rect 33048 8041 33057 8075
rect 33057 8041 33091 8075
rect 33091 8041 33100 8075
rect 33048 8032 33100 8041
rect 33508 8032 33560 8084
rect 40592 8032 40644 8084
rect 42248 8075 42300 8084
rect 42248 8041 42257 8075
rect 42257 8041 42291 8075
rect 42291 8041 42300 8075
rect 42248 8032 42300 8041
rect 50160 8075 50212 8084
rect 50160 8041 50169 8075
rect 50169 8041 50203 8075
rect 50203 8041 50212 8075
rect 50160 8032 50212 8041
rect 53288 8032 53340 8084
rect 49516 7964 49568 8016
rect 50712 7964 50764 8016
rect 16672 7828 16724 7880
rect 17132 7828 17184 7880
rect 16120 7760 16172 7812
rect 16212 7760 16264 7812
rect 17316 7760 17368 7812
rect 6644 7692 6696 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 11060 7735 11112 7744
rect 6920 7692 6972 7701
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 11520 7692 11572 7744
rect 17776 7692 17828 7744
rect 19340 7828 19392 7880
rect 20812 7760 20864 7812
rect 22744 7828 22796 7880
rect 27528 7896 27580 7948
rect 27804 7896 27856 7948
rect 33600 7939 33652 7948
rect 26884 7871 26936 7880
rect 22192 7760 22244 7812
rect 25136 7760 25188 7812
rect 26884 7837 26893 7871
rect 26893 7837 26927 7871
rect 26927 7837 26936 7871
rect 26884 7828 26936 7837
rect 27160 7871 27212 7880
rect 27160 7837 27169 7871
rect 27169 7837 27203 7871
rect 27203 7837 27212 7871
rect 27160 7828 27212 7837
rect 28172 7828 28224 7880
rect 28632 7871 28684 7880
rect 28632 7837 28641 7871
rect 28641 7837 28675 7871
rect 28675 7837 28684 7871
rect 28632 7828 28684 7837
rect 33600 7905 33609 7939
rect 33609 7905 33643 7939
rect 33643 7905 33652 7939
rect 33600 7896 33652 7905
rect 39120 7896 39172 7948
rect 40040 7896 40092 7948
rect 40684 7896 40736 7948
rect 42708 7896 42760 7948
rect 50620 7939 50672 7948
rect 50620 7905 50629 7939
rect 50629 7905 50663 7939
rect 50663 7905 50672 7939
rect 50620 7896 50672 7905
rect 52644 7939 52696 7948
rect 52644 7905 52653 7939
rect 52653 7905 52687 7939
rect 52687 7905 52696 7939
rect 52644 7896 52696 7905
rect 30472 7828 30524 7880
rect 36176 7828 36228 7880
rect 36360 7828 36412 7880
rect 38384 7828 38436 7880
rect 50252 7828 50304 7880
rect 29552 7760 29604 7812
rect 33232 7760 33284 7812
rect 42616 7803 42668 7812
rect 42616 7769 42625 7803
rect 42625 7769 42659 7803
rect 42659 7769 42668 7803
rect 42616 7760 42668 7769
rect 45192 7760 45244 7812
rect 53104 7760 53156 7812
rect 20996 7735 21048 7744
rect 20996 7701 21005 7735
rect 21005 7701 21039 7735
rect 21039 7701 21048 7735
rect 20996 7692 21048 7701
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 23848 7692 23900 7744
rect 26700 7735 26752 7744
rect 26700 7701 26709 7735
rect 26709 7701 26743 7735
rect 26743 7701 26752 7735
rect 26700 7692 26752 7701
rect 27068 7735 27120 7744
rect 27068 7701 27077 7735
rect 27077 7701 27111 7735
rect 27111 7701 27120 7735
rect 27068 7692 27120 7701
rect 27804 7735 27856 7744
rect 27804 7701 27813 7735
rect 27813 7701 27847 7735
rect 27847 7701 27856 7735
rect 27804 7692 27856 7701
rect 28172 7735 28224 7744
rect 28172 7701 28181 7735
rect 28181 7701 28215 7735
rect 28215 7701 28224 7735
rect 28172 7692 28224 7701
rect 34336 7692 34388 7744
rect 42800 7692 42852 7744
rect 43904 7692 43956 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 12716 7488 12768 7540
rect 13176 7488 13228 7540
rect 16856 7488 16908 7540
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 6920 7420 6972 7472
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6644 7395 6696 7404
rect 6644 7361 6678 7395
rect 6678 7361 6696 7395
rect 6644 7352 6696 7361
rect 3240 7216 3292 7268
rect 9680 7395 9732 7404
rect 9680 7361 9714 7395
rect 9714 7361 9732 7395
rect 13912 7395 13964 7404
rect 9680 7352 9732 7361
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 14280 7420 14332 7472
rect 19248 7420 19300 7472
rect 14464 7352 14516 7404
rect 15200 7352 15252 7404
rect 6092 7148 6144 7200
rect 6368 7148 6420 7200
rect 14648 7284 14700 7336
rect 11428 7216 11480 7268
rect 14096 7216 14148 7268
rect 17132 7395 17184 7404
rect 17132 7361 17146 7395
rect 17146 7361 17180 7395
rect 17180 7361 17184 7395
rect 17132 7352 17184 7361
rect 17684 7352 17736 7404
rect 19892 7284 19944 7336
rect 20628 7395 20680 7404
rect 20628 7361 20637 7395
rect 20637 7361 20671 7395
rect 20671 7361 20680 7395
rect 20628 7352 20680 7361
rect 20720 7284 20772 7336
rect 21824 7284 21876 7336
rect 16120 7216 16172 7268
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 22744 7395 22796 7404
rect 22744 7361 22753 7395
rect 22753 7361 22787 7395
rect 22787 7361 22796 7395
rect 22744 7352 22796 7361
rect 23756 7420 23808 7472
rect 26700 7420 26752 7472
rect 27712 7420 27764 7472
rect 28632 7420 28684 7472
rect 32864 7420 32916 7472
rect 36360 7488 36412 7540
rect 36544 7488 36596 7540
rect 37004 7488 37056 7540
rect 53104 7531 53156 7540
rect 53104 7497 53113 7531
rect 53113 7497 53147 7531
rect 53147 7497 53156 7531
rect 53104 7488 53156 7497
rect 36452 7420 36504 7472
rect 37096 7420 37148 7472
rect 37464 7420 37516 7472
rect 40684 7420 40736 7472
rect 52920 7420 52972 7472
rect 28172 7352 28224 7404
rect 32312 7395 32364 7404
rect 32312 7361 32321 7395
rect 32321 7361 32355 7395
rect 32355 7361 32364 7395
rect 32312 7352 32364 7361
rect 32404 7395 32456 7404
rect 32404 7361 32413 7395
rect 32413 7361 32447 7395
rect 32447 7361 32456 7395
rect 32404 7352 32456 7361
rect 9588 7148 9640 7200
rect 12532 7148 12584 7200
rect 21916 7148 21968 7200
rect 23480 7284 23532 7336
rect 26792 7284 26844 7336
rect 30932 7284 30984 7336
rect 32496 7284 32548 7336
rect 33140 7352 33192 7404
rect 35440 7352 35492 7404
rect 38384 7352 38436 7404
rect 43720 7395 43772 7404
rect 43720 7361 43729 7395
rect 43729 7361 43763 7395
rect 43763 7361 43772 7395
rect 43720 7352 43772 7361
rect 44548 7352 44600 7404
rect 45284 7352 45336 7404
rect 47308 7352 47360 7404
rect 53012 7395 53064 7404
rect 53012 7361 53021 7395
rect 53021 7361 53055 7395
rect 53055 7361 53064 7395
rect 53012 7352 53064 7361
rect 46940 7284 46992 7336
rect 22928 7148 22980 7200
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 27988 7148 28040 7200
rect 32128 7191 32180 7200
rect 32128 7157 32137 7191
rect 32137 7157 32171 7191
rect 32171 7157 32180 7191
rect 32128 7148 32180 7157
rect 32404 7148 32456 7200
rect 33324 7148 33376 7200
rect 35348 7216 35400 7268
rect 37004 7216 37056 7268
rect 42708 7216 42760 7268
rect 35992 7191 36044 7200
rect 35992 7157 36001 7191
rect 36001 7157 36035 7191
rect 36035 7157 36044 7191
rect 35992 7148 36044 7157
rect 36176 7191 36228 7200
rect 36176 7157 36185 7191
rect 36185 7157 36219 7191
rect 36219 7157 36228 7191
rect 36176 7148 36228 7157
rect 37832 7191 37884 7200
rect 37832 7157 37841 7191
rect 37841 7157 37875 7191
rect 37875 7157 37884 7191
rect 37832 7148 37884 7157
rect 45192 7148 45244 7200
rect 46204 7191 46256 7200
rect 46204 7157 46213 7191
rect 46213 7157 46247 7191
rect 46247 7157 46256 7191
rect 46204 7148 46256 7157
rect 46572 7191 46624 7200
rect 46572 7157 46581 7191
rect 46581 7157 46615 7191
rect 46615 7157 46624 7191
rect 46572 7148 46624 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9680 6944 9732 6996
rect 13268 6944 13320 6996
rect 13728 6944 13780 6996
rect 14648 6944 14700 6996
rect 16120 6944 16172 6996
rect 2044 6876 2096 6928
rect 3792 6876 3844 6928
rect 8024 6876 8076 6928
rect 9956 6876 10008 6928
rect 16212 6876 16264 6928
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2780 6740 2832 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 9680 6808 9732 6860
rect 7104 6740 7156 6792
rect 7472 6740 7524 6792
rect 11060 6740 11112 6792
rect 13084 6783 13136 6792
rect 13084 6749 13091 6783
rect 13091 6749 13136 6783
rect 13084 6740 13136 6749
rect 7840 6672 7892 6724
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7104 6604 7156 6656
rect 9956 6604 10008 6656
rect 13728 6740 13780 6792
rect 14096 6783 14148 6792
rect 14096 6749 14112 6783
rect 14112 6749 14146 6783
rect 14146 6749 14148 6783
rect 14096 6740 14148 6749
rect 14280 6740 14332 6792
rect 14924 6808 14976 6860
rect 14648 6740 14700 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 13268 6715 13320 6724
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 16856 6876 16908 6928
rect 16672 6740 16724 6792
rect 13268 6672 13320 6681
rect 14188 6604 14240 6656
rect 19432 6944 19484 6996
rect 21548 6987 21600 6996
rect 21548 6953 21557 6987
rect 21557 6953 21591 6987
rect 21591 6953 21600 6987
rect 21548 6944 21600 6953
rect 21640 6944 21692 6996
rect 25136 6944 25188 6996
rect 32312 6944 32364 6996
rect 35992 6987 36044 6996
rect 35992 6953 36001 6987
rect 36001 6953 36035 6987
rect 36035 6953 36044 6987
rect 35992 6944 36044 6953
rect 36176 6944 36228 6996
rect 46572 6944 46624 6996
rect 20996 6919 21048 6928
rect 20996 6885 21005 6919
rect 21005 6885 21039 6919
rect 21039 6885 21048 6919
rect 20996 6876 21048 6885
rect 17316 6783 17368 6792
rect 17316 6749 17326 6783
rect 17326 6749 17360 6783
rect 17360 6749 17368 6783
rect 17316 6740 17368 6749
rect 17684 6783 17736 6792
rect 17684 6749 17698 6783
rect 17698 6749 17732 6783
rect 17732 6749 17736 6783
rect 17684 6740 17736 6749
rect 19892 6740 19944 6792
rect 20076 6672 20128 6724
rect 20260 6740 20312 6792
rect 21916 6808 21968 6860
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 26056 6808 26108 6860
rect 30932 6808 30984 6860
rect 37004 6876 37056 6928
rect 37372 6876 37424 6928
rect 37556 6808 37608 6860
rect 38476 6808 38528 6860
rect 41880 6919 41932 6928
rect 41880 6885 41889 6919
rect 41889 6885 41923 6919
rect 41923 6885 41932 6919
rect 41880 6876 41932 6885
rect 22284 6783 22336 6792
rect 22284 6749 22293 6783
rect 22293 6749 22327 6783
rect 22327 6749 22336 6783
rect 22284 6740 22336 6749
rect 22376 6740 22428 6792
rect 20628 6672 20680 6724
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 16672 6604 16724 6656
rect 16948 6604 17000 6656
rect 17868 6647 17920 6656
rect 17868 6613 17877 6647
rect 17877 6613 17911 6647
rect 17911 6613 17920 6647
rect 17868 6604 17920 6613
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 22468 6672 22520 6724
rect 29552 6740 29604 6792
rect 31024 6783 31076 6792
rect 31024 6749 31033 6783
rect 31033 6749 31067 6783
rect 31067 6749 31076 6783
rect 31024 6740 31076 6749
rect 32128 6672 32180 6724
rect 33140 6672 33192 6724
rect 20536 6604 20588 6613
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 21272 6604 21324 6613
rect 26240 6604 26292 6656
rect 31392 6604 31444 6656
rect 32404 6647 32456 6656
rect 32404 6613 32413 6647
rect 32413 6613 32447 6647
rect 32447 6613 32456 6647
rect 33232 6647 33284 6656
rect 32404 6604 32456 6613
rect 33232 6613 33241 6647
rect 33241 6613 33275 6647
rect 33275 6613 33284 6647
rect 33232 6604 33284 6613
rect 33324 6647 33376 6656
rect 33324 6613 33333 6647
rect 33333 6613 33367 6647
rect 33367 6613 33376 6647
rect 34152 6672 34204 6724
rect 35440 6672 35492 6724
rect 37004 6740 37056 6792
rect 37280 6783 37332 6792
rect 37280 6749 37289 6783
rect 37289 6749 37323 6783
rect 37323 6749 37332 6783
rect 37280 6740 37332 6749
rect 38384 6740 38436 6792
rect 40132 6740 40184 6792
rect 40408 6783 40460 6792
rect 40408 6749 40417 6783
rect 40417 6749 40451 6783
rect 40451 6749 40460 6783
rect 40408 6740 40460 6749
rect 40960 6740 41012 6792
rect 42892 6851 42944 6860
rect 42892 6817 42901 6851
rect 42901 6817 42935 6851
rect 42935 6817 42944 6851
rect 42892 6808 42944 6817
rect 43168 6808 43220 6860
rect 41696 6783 41748 6792
rect 41696 6749 41705 6783
rect 41705 6749 41739 6783
rect 41739 6749 41748 6783
rect 41696 6740 41748 6749
rect 35992 6715 36044 6724
rect 35992 6681 36017 6715
rect 36017 6681 36044 6715
rect 35992 6672 36044 6681
rect 33324 6604 33376 6613
rect 35348 6604 35400 6656
rect 38292 6604 38344 6656
rect 40224 6604 40276 6656
rect 41052 6672 41104 6724
rect 40868 6604 40920 6656
rect 40960 6604 41012 6656
rect 41972 6740 42024 6792
rect 42984 6740 43036 6792
rect 43076 6740 43128 6792
rect 45560 6740 45612 6792
rect 46572 6783 46624 6792
rect 43352 6672 43404 6724
rect 43720 6672 43772 6724
rect 46572 6749 46581 6783
rect 46581 6749 46615 6783
rect 46615 6749 46624 6783
rect 46572 6740 46624 6749
rect 49148 6783 49200 6792
rect 49148 6749 49157 6783
rect 49157 6749 49191 6783
rect 49191 6749 49200 6783
rect 49148 6740 49200 6749
rect 50620 6740 50672 6792
rect 46204 6672 46256 6724
rect 47952 6647 48004 6656
rect 47952 6613 47961 6647
rect 47961 6613 47995 6647
rect 47995 6613 48004 6647
rect 47952 6604 48004 6613
rect 49332 6672 49384 6724
rect 49148 6604 49200 6656
rect 49424 6604 49476 6656
rect 52644 6647 52696 6656
rect 52644 6613 52653 6647
rect 52653 6613 52687 6647
rect 52687 6613 52696 6647
rect 52644 6604 52696 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 10876 6332 10928 6384
rect 15292 6400 15344 6452
rect 17316 6400 17368 6452
rect 20168 6400 20220 6452
rect 25780 6400 25832 6452
rect 30012 6400 30064 6452
rect 19984 6332 20036 6384
rect 2964 6264 3016 6316
rect 5172 6264 5224 6316
rect 9864 6307 9916 6316
rect 9864 6273 9898 6307
rect 9898 6273 9916 6307
rect 9864 6264 9916 6273
rect 10600 6264 10652 6316
rect 13268 6264 13320 6316
rect 16212 6264 16264 6316
rect 19432 6264 19484 6316
rect 20536 6264 20588 6316
rect 21456 6264 21508 6316
rect 24400 6332 24452 6384
rect 22836 6264 22888 6316
rect 25872 6264 25924 6316
rect 26056 6307 26108 6316
rect 26056 6273 26065 6307
rect 26065 6273 26099 6307
rect 26099 6273 26108 6307
rect 26056 6264 26108 6273
rect 26240 6307 26292 6316
rect 26240 6273 26249 6307
rect 26249 6273 26283 6307
rect 26283 6273 26292 6307
rect 26240 6264 26292 6273
rect 26792 6264 26844 6316
rect 29092 6264 29144 6316
rect 2596 6196 2648 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 11888 6196 11940 6248
rect 20812 6196 20864 6248
rect 22100 6239 22152 6248
rect 22100 6205 22109 6239
rect 22109 6205 22143 6239
rect 22143 6205 22152 6239
rect 22284 6239 22336 6248
rect 22100 6196 22152 6205
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22468 6196 22520 6248
rect 29736 6307 29788 6316
rect 29736 6273 29745 6307
rect 29745 6273 29779 6307
rect 29779 6273 29788 6307
rect 29736 6264 29788 6273
rect 31116 6400 31168 6452
rect 30656 6332 30708 6384
rect 30932 6332 30984 6384
rect 33324 6400 33376 6452
rect 32220 6332 32272 6384
rect 36084 6400 36136 6452
rect 36268 6400 36320 6452
rect 30472 6307 30524 6316
rect 30472 6273 30481 6307
rect 30481 6273 30515 6307
rect 30515 6273 30524 6307
rect 30472 6264 30524 6273
rect 31024 6264 31076 6316
rect 33416 6264 33468 6316
rect 34152 6307 34204 6316
rect 34152 6273 34161 6307
rect 34161 6273 34195 6307
rect 34195 6273 34204 6307
rect 34152 6264 34204 6273
rect 34244 6307 34296 6316
rect 34244 6273 34253 6307
rect 34253 6273 34287 6307
rect 34287 6273 34296 6307
rect 37740 6332 37792 6384
rect 38568 6332 38620 6384
rect 40408 6400 40460 6452
rect 46940 6443 46992 6452
rect 46940 6409 46949 6443
rect 46949 6409 46983 6443
rect 46983 6409 46992 6443
rect 46940 6400 46992 6409
rect 47032 6400 47084 6452
rect 48872 6400 48924 6452
rect 34244 6264 34296 6273
rect 35348 6264 35400 6316
rect 8300 6128 8352 6180
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 8852 6060 8904 6112
rect 14280 6060 14332 6112
rect 19984 6060 20036 6112
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 20720 6128 20772 6180
rect 21640 6060 21692 6112
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 22192 6128 22244 6180
rect 34796 6196 34848 6248
rect 35992 6196 36044 6248
rect 36360 6264 36412 6316
rect 36912 6264 36964 6316
rect 39396 6307 39448 6316
rect 39396 6273 39405 6307
rect 39405 6273 39439 6307
rect 39439 6273 39448 6307
rect 39396 6264 39448 6273
rect 40132 6332 40184 6384
rect 22468 6060 22520 6112
rect 25596 6060 25648 6112
rect 26148 6060 26200 6112
rect 33692 6128 33744 6180
rect 40868 6196 40920 6248
rect 41880 6264 41932 6316
rect 43076 6264 43128 6316
rect 43536 6264 43588 6316
rect 46572 6307 46624 6316
rect 46572 6273 46581 6307
rect 46581 6273 46615 6307
rect 46615 6273 46624 6307
rect 46572 6264 46624 6273
rect 46664 6307 46716 6316
rect 46664 6273 46673 6307
rect 46673 6273 46707 6307
rect 46707 6273 46716 6307
rect 46664 6264 46716 6273
rect 47124 6264 47176 6316
rect 47308 6264 47360 6316
rect 41604 6196 41656 6248
rect 43260 6239 43312 6248
rect 43260 6205 43269 6239
rect 43269 6205 43303 6239
rect 43303 6205 43312 6239
rect 43260 6196 43312 6205
rect 29644 6060 29696 6112
rect 34428 6103 34480 6112
rect 34428 6069 34437 6103
rect 34437 6069 34471 6103
rect 34471 6069 34480 6103
rect 34428 6060 34480 6069
rect 34704 6060 34756 6112
rect 38568 6128 38620 6180
rect 39396 6128 39448 6180
rect 42708 6128 42760 6180
rect 43720 6196 43772 6248
rect 48044 6239 48096 6248
rect 48044 6205 48053 6239
rect 48053 6205 48087 6239
rect 48087 6205 48096 6239
rect 48044 6196 48096 6205
rect 36728 6060 36780 6112
rect 39212 6103 39264 6112
rect 39212 6069 39221 6103
rect 39221 6069 39255 6103
rect 39255 6069 39264 6103
rect 39212 6060 39264 6069
rect 41512 6060 41564 6112
rect 41696 6060 41748 6112
rect 45560 6060 45612 6112
rect 46756 6060 46808 6112
rect 46848 6060 46900 6112
rect 48596 6060 48648 6112
rect 49424 6060 49476 6112
rect 50160 6103 50212 6112
rect 50160 6069 50169 6103
rect 50169 6069 50203 6103
rect 50203 6069 50212 6103
rect 50160 6060 50212 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 7840 5899 7892 5908
rect 7840 5865 7849 5899
rect 7849 5865 7883 5899
rect 7883 5865 7892 5899
rect 7840 5856 7892 5865
rect 9864 5856 9916 5908
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 20628 5856 20680 5908
rect 22192 5856 22244 5908
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 2596 5763 2648 5772
rect 2596 5729 2605 5763
rect 2605 5729 2639 5763
rect 2639 5729 2648 5763
rect 2596 5720 2648 5729
rect 3608 5720 3660 5772
rect 12440 5788 12492 5840
rect 13084 5788 13136 5840
rect 19892 5788 19944 5840
rect 21456 5831 21508 5840
rect 21456 5797 21465 5831
rect 21465 5797 21499 5831
rect 21499 5797 21508 5831
rect 21456 5788 21508 5797
rect 22100 5788 22152 5840
rect 11060 5720 11112 5772
rect 20628 5720 20680 5772
rect 21732 5720 21784 5772
rect 41880 5856 41932 5908
rect 27620 5831 27672 5840
rect 27620 5797 27629 5831
rect 27629 5797 27663 5831
rect 27663 5797 27672 5831
rect 27620 5788 27672 5797
rect 30932 5831 30984 5840
rect 30932 5797 30941 5831
rect 30941 5797 30975 5831
rect 30975 5797 30984 5831
rect 30932 5788 30984 5797
rect 23480 5720 23532 5772
rect 24124 5720 24176 5772
rect 3148 5652 3200 5704
rect 6092 5652 6144 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10324 5652 10376 5704
rect 13820 5652 13872 5704
rect 14464 5695 14516 5704
rect 4252 5584 4304 5636
rect 7932 5584 7984 5636
rect 9496 5584 9548 5636
rect 12900 5584 12952 5636
rect 3332 5516 3384 5568
rect 3608 5516 3660 5568
rect 5172 5516 5224 5568
rect 7196 5516 7248 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 16396 5652 16448 5704
rect 19984 5652 20036 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 21916 5695 21968 5704
rect 21916 5661 21925 5695
rect 21925 5661 21959 5695
rect 21959 5661 21968 5695
rect 21916 5652 21968 5661
rect 29092 5720 29144 5772
rect 29552 5763 29604 5772
rect 29552 5729 29561 5763
rect 29561 5729 29595 5763
rect 29595 5729 29604 5763
rect 29552 5720 29604 5729
rect 19432 5584 19484 5636
rect 21180 5516 21232 5568
rect 26792 5652 26844 5704
rect 29644 5652 29696 5704
rect 24860 5584 24912 5636
rect 26332 5584 26384 5636
rect 26976 5584 27028 5636
rect 32220 5720 32272 5772
rect 33048 5788 33100 5840
rect 34704 5788 34756 5840
rect 35532 5788 35584 5840
rect 47308 5856 47360 5908
rect 47492 5856 47544 5908
rect 43352 5831 43404 5840
rect 43352 5797 43361 5831
rect 43361 5797 43395 5831
rect 43395 5797 43404 5831
rect 43352 5788 43404 5797
rect 34704 5695 34756 5704
rect 34704 5661 34713 5695
rect 34713 5661 34747 5695
rect 34747 5661 34756 5695
rect 34704 5652 34756 5661
rect 33140 5584 33192 5636
rect 25872 5516 25924 5568
rect 26056 5516 26108 5568
rect 32496 5516 32548 5568
rect 36360 5652 36412 5704
rect 38200 5652 38252 5704
rect 41236 5652 41288 5704
rect 41512 5695 41564 5704
rect 41512 5661 41521 5695
rect 41521 5661 41555 5695
rect 41555 5661 41564 5695
rect 41512 5652 41564 5661
rect 41972 5695 42024 5704
rect 41972 5661 41981 5695
rect 41981 5661 42015 5695
rect 42015 5661 42024 5695
rect 41972 5652 42024 5661
rect 43260 5720 43312 5772
rect 47032 5788 47084 5840
rect 48044 5788 48096 5840
rect 46572 5720 46624 5772
rect 45100 5695 45152 5704
rect 45100 5661 45109 5695
rect 45109 5661 45143 5695
rect 45143 5661 45152 5695
rect 45100 5652 45152 5661
rect 46664 5652 46716 5704
rect 35164 5584 35216 5636
rect 35900 5627 35952 5636
rect 35440 5516 35492 5568
rect 35900 5593 35909 5627
rect 35909 5593 35943 5627
rect 35943 5593 35952 5627
rect 35900 5584 35952 5593
rect 36728 5584 36780 5636
rect 40224 5584 40276 5636
rect 40408 5584 40460 5636
rect 40868 5584 40920 5636
rect 40960 5516 41012 5568
rect 45652 5584 45704 5636
rect 41972 5516 42024 5568
rect 43720 5516 43772 5568
rect 45284 5559 45336 5568
rect 45284 5525 45293 5559
rect 45293 5525 45327 5559
rect 45327 5525 45336 5559
rect 45284 5516 45336 5525
rect 47124 5720 47176 5772
rect 47400 5652 47452 5704
rect 49148 5652 49200 5704
rect 50620 5856 50672 5908
rect 47032 5627 47084 5636
rect 47032 5593 47041 5627
rect 47041 5593 47075 5627
rect 47075 5593 47084 5627
rect 47032 5584 47084 5593
rect 48780 5627 48832 5636
rect 47952 5516 48004 5568
rect 48780 5593 48789 5627
rect 48789 5593 48823 5627
rect 48823 5593 48832 5627
rect 48780 5584 48832 5593
rect 50160 5516 50212 5568
rect 51080 5516 51132 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 1676 5312 1728 5364
rect 7104 5312 7156 5364
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 8300 5312 8352 5364
rect 14464 5312 14516 5364
rect 17776 5312 17828 5364
rect 20812 5312 20864 5364
rect 21272 5355 21324 5364
rect 21272 5321 21281 5355
rect 21281 5321 21315 5355
rect 21315 5321 21324 5355
rect 21272 5312 21324 5321
rect 24860 5355 24912 5364
rect 24860 5321 24869 5355
rect 24869 5321 24903 5355
rect 24903 5321 24912 5355
rect 24860 5312 24912 5321
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 1860 5287 1912 5296
rect 1860 5253 1869 5287
rect 1869 5253 1903 5287
rect 1903 5253 1912 5287
rect 1860 5244 1912 5253
rect 10048 5244 10100 5296
rect 10324 5244 10376 5296
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 4988 5176 5040 5228
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 7104 5219 7156 5228
rect 6920 5176 6972 5185
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 14096 5244 14148 5296
rect 21824 5244 21876 5296
rect 33048 5244 33100 5296
rect 15384 5176 15436 5228
rect 16764 5176 16816 5228
rect 19340 5176 19392 5228
rect 20536 5176 20588 5228
rect 24216 5219 24268 5228
rect 24216 5185 24225 5219
rect 24225 5185 24259 5219
rect 24259 5185 24268 5219
rect 24216 5176 24268 5185
rect 25596 5219 25648 5228
rect 25596 5185 25605 5219
rect 25605 5185 25639 5219
rect 25639 5185 25648 5219
rect 25596 5176 25648 5185
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 25964 5219 26016 5228
rect 25964 5185 25973 5219
rect 25973 5185 26007 5219
rect 26007 5185 26016 5219
rect 25964 5176 26016 5185
rect 26148 5219 26200 5228
rect 26148 5185 26157 5219
rect 26157 5185 26191 5219
rect 26191 5185 26200 5219
rect 26148 5176 26200 5185
rect 27620 5176 27672 5228
rect 34428 5312 34480 5364
rect 35348 5244 35400 5296
rect 35992 5312 36044 5364
rect 36084 5312 36136 5364
rect 40316 5312 40368 5364
rect 39212 5244 39264 5296
rect 40224 5244 40276 5296
rect 41052 5244 41104 5296
rect 51080 5287 51132 5296
rect 51080 5253 51114 5287
rect 51114 5253 51132 5287
rect 51080 5244 51132 5253
rect 2780 5040 2832 5092
rect 9588 5040 9640 5092
rect 10140 5040 10192 5092
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 3884 4972 3936 5024
rect 5264 4972 5316 5024
rect 6736 4972 6788 5024
rect 10416 4972 10468 5024
rect 15476 4972 15528 5024
rect 22468 5108 22520 5160
rect 24492 5108 24544 5160
rect 25872 5151 25924 5160
rect 25872 5117 25881 5151
rect 25881 5117 25915 5151
rect 25915 5117 25924 5151
rect 25872 5108 25924 5117
rect 24768 5040 24820 5092
rect 33048 5108 33100 5160
rect 34336 5176 34388 5228
rect 48596 5176 48648 5228
rect 37924 5108 37976 5160
rect 30472 4972 30524 5024
rect 35256 5040 35308 5092
rect 33508 4972 33560 5024
rect 34244 4972 34296 5024
rect 35900 4972 35952 5024
rect 41972 5040 42024 5092
rect 40132 4972 40184 5024
rect 48964 4972 49016 5024
rect 52184 5015 52236 5024
rect 52184 4981 52193 5015
rect 52193 4981 52227 5015
rect 52227 4981 52236 5015
rect 52184 4972 52236 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 7472 4811 7524 4820
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 5172 4743 5224 4752
rect 5172 4709 5181 4743
rect 5181 4709 5215 4743
rect 5215 4709 5224 4743
rect 5172 4700 5224 4709
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 10048 4768 10100 4820
rect 16764 4768 16816 4820
rect 24216 4768 24268 4820
rect 30656 4811 30708 4820
rect 30656 4777 30665 4811
rect 30665 4777 30699 4811
rect 30699 4777 30708 4811
rect 30656 4768 30708 4777
rect 35532 4768 35584 4820
rect 35992 4811 36044 4820
rect 35992 4777 36001 4811
rect 36001 4777 36035 4811
rect 36035 4777 36044 4811
rect 35992 4768 36044 4777
rect 38660 4768 38712 4820
rect 48780 4768 48832 4820
rect 9588 4700 9640 4752
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3884 4564 3936 4616
rect 5540 4564 5592 4616
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 3700 4496 3752 4548
rect 6920 4564 6972 4616
rect 7748 4564 7800 4616
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 9772 4564 9824 4616
rect 10416 4607 10468 4616
rect 10416 4573 10450 4607
rect 10450 4573 10468 4607
rect 10416 4564 10468 4573
rect 13636 4564 13688 4616
rect 19524 4700 19576 4752
rect 16396 4632 16448 4684
rect 6644 4496 6696 4548
rect 13544 4496 13596 4548
rect 1584 4428 1636 4480
rect 2964 4428 3016 4480
rect 5172 4428 5224 4480
rect 7104 4428 7156 4480
rect 7840 4428 7892 4480
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 15752 4428 15804 4437
rect 16580 4496 16632 4548
rect 17776 4496 17828 4548
rect 22284 4632 22336 4684
rect 23296 4632 23348 4684
rect 26056 4700 26108 4752
rect 29000 4700 29052 4752
rect 33232 4700 33284 4752
rect 33876 4700 33928 4752
rect 20260 4564 20312 4616
rect 22652 4564 22704 4616
rect 24492 4607 24544 4616
rect 24492 4573 24502 4607
rect 24502 4573 24536 4607
rect 24536 4573 24544 4607
rect 24492 4564 24544 4573
rect 24860 4607 24912 4616
rect 24860 4573 24874 4607
rect 24874 4573 24908 4607
rect 24908 4573 24912 4607
rect 24860 4564 24912 4573
rect 25136 4564 25188 4616
rect 26148 4564 26200 4616
rect 34244 4632 34296 4684
rect 37464 4700 37516 4752
rect 40316 4700 40368 4752
rect 48872 4700 48924 4752
rect 36084 4632 36136 4684
rect 39764 4632 39816 4684
rect 40040 4632 40092 4684
rect 29552 4564 29604 4616
rect 30472 4607 30524 4616
rect 30472 4573 30481 4607
rect 30481 4573 30515 4607
rect 30515 4573 30524 4607
rect 30472 4564 30524 4573
rect 31116 4607 31168 4616
rect 31116 4573 31125 4607
rect 31125 4573 31159 4607
rect 31159 4573 31168 4607
rect 31116 4564 31168 4573
rect 31576 4564 31628 4616
rect 33324 4607 33376 4616
rect 33324 4573 33333 4607
rect 33333 4573 33367 4607
rect 33367 4573 33376 4607
rect 33324 4564 33376 4573
rect 33508 4607 33560 4616
rect 33508 4573 33517 4607
rect 33517 4573 33551 4607
rect 33551 4573 33560 4607
rect 33508 4564 33560 4573
rect 33692 4607 33744 4616
rect 33692 4573 33701 4607
rect 33701 4573 33735 4607
rect 33735 4573 33744 4607
rect 33692 4564 33744 4573
rect 35256 4585 35308 4616
rect 35256 4564 35265 4585
rect 35265 4564 35299 4585
rect 35299 4564 35308 4585
rect 35440 4607 35492 4616
rect 35440 4573 35455 4607
rect 35455 4573 35492 4607
rect 35440 4564 35492 4573
rect 35716 4564 35768 4616
rect 35900 4564 35952 4616
rect 37556 4564 37608 4616
rect 39856 4607 39908 4616
rect 39856 4573 39865 4607
rect 39865 4573 39899 4607
rect 39899 4573 39908 4607
rect 39856 4564 39908 4573
rect 40132 4607 40184 4616
rect 40132 4573 40141 4607
rect 40141 4573 40175 4607
rect 40175 4573 40184 4607
rect 40132 4564 40184 4573
rect 40776 4632 40828 4684
rect 45468 4632 45520 4684
rect 46296 4632 46348 4684
rect 47124 4675 47176 4684
rect 47124 4641 47133 4675
rect 47133 4641 47167 4675
rect 47167 4641 47176 4675
rect 47124 4632 47176 4641
rect 47492 4632 47544 4684
rect 48044 4632 48096 4684
rect 48688 4607 48740 4616
rect 48688 4573 48697 4607
rect 48697 4573 48731 4607
rect 48731 4573 48740 4607
rect 48688 4564 48740 4573
rect 48872 4607 48924 4616
rect 48872 4573 48881 4607
rect 48881 4573 48915 4607
rect 48915 4573 48924 4607
rect 48872 4564 48924 4573
rect 49148 4564 49200 4616
rect 19524 4539 19576 4548
rect 19524 4505 19533 4539
rect 19533 4505 19567 4539
rect 19567 4505 19576 4539
rect 19524 4496 19576 4505
rect 20444 4496 20496 4548
rect 24308 4496 24360 4548
rect 25872 4496 25924 4548
rect 27988 4539 28040 4548
rect 27988 4505 27997 4539
rect 27997 4505 28031 4539
rect 28031 4505 28040 4539
rect 27988 4496 28040 4505
rect 30196 4496 30248 4548
rect 30932 4496 30984 4548
rect 31300 4539 31352 4548
rect 31300 4505 31309 4539
rect 31309 4505 31343 4539
rect 31343 4505 31352 4539
rect 31300 4496 31352 4505
rect 33140 4496 33192 4548
rect 33600 4539 33652 4548
rect 33600 4505 33609 4539
rect 33609 4505 33643 4539
rect 33643 4505 33652 4539
rect 33600 4496 33652 4505
rect 19432 4428 19484 4480
rect 22100 4428 22152 4480
rect 27712 4428 27764 4480
rect 31576 4428 31628 4480
rect 40316 4496 40368 4548
rect 45100 4496 45152 4548
rect 48320 4496 48372 4548
rect 48964 4539 49016 4548
rect 48964 4505 48973 4539
rect 48973 4505 49007 4539
rect 49007 4505 49016 4539
rect 48964 4496 49016 4505
rect 33968 4428 34020 4480
rect 34244 4428 34296 4480
rect 37556 4428 37608 4480
rect 37740 4428 37792 4480
rect 41236 4428 41288 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 6644 4267 6696 4276
rect 2780 4088 2832 4140
rect 3884 4156 3936 4208
rect 4160 4156 4212 4208
rect 4988 4156 5040 4208
rect 5080 4156 5132 4208
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 6736 4267 6788 4276
rect 6736 4233 6745 4267
rect 6745 4233 6779 4267
rect 6779 4233 6788 4267
rect 7932 4267 7984 4276
rect 6736 4224 6788 4233
rect 7932 4233 7941 4267
rect 7941 4233 7975 4267
rect 7975 4233 7984 4267
rect 7932 4224 7984 4233
rect 3700 4088 3752 4140
rect 5448 4156 5500 4208
rect 5540 4088 5592 4140
rect 6552 4088 6604 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 9312 4156 9364 4208
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2964 4020 3016 4072
rect 6644 4020 6696 4072
rect 6736 4020 6788 4072
rect 8392 4088 8444 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10416 4088 10468 4140
rect 12532 4156 12584 4208
rect 13820 4156 13872 4208
rect 12992 4088 13044 4140
rect 8024 4020 8076 4072
rect 20168 4224 20220 4276
rect 24492 4224 24544 4276
rect 15016 4156 15068 4208
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 16212 4088 16264 4140
rect 24860 4156 24912 4208
rect 25780 4224 25832 4276
rect 31300 4224 31352 4276
rect 33048 4224 33100 4276
rect 37464 4224 37516 4276
rect 41052 4224 41104 4276
rect 43812 4267 43864 4276
rect 19064 4088 19116 4140
rect 19432 4088 19484 4140
rect 23296 4088 23348 4140
rect 23572 4088 23624 4140
rect 24400 4088 24452 4140
rect 25504 4088 25556 4140
rect 25872 4088 25924 4140
rect 29092 4156 29144 4208
rect 22376 4020 22428 4072
rect 22468 4063 22520 4072
rect 22468 4029 22477 4063
rect 22477 4029 22511 4063
rect 22511 4029 22520 4063
rect 22468 4020 22520 4029
rect 23020 4020 23072 4072
rect 3240 3952 3292 4004
rect 2136 3884 2188 3936
rect 5080 3952 5132 4004
rect 6736 3884 6788 3936
rect 8024 3884 8076 3936
rect 8116 3884 8168 3936
rect 10140 3952 10192 4004
rect 10600 3952 10652 4004
rect 10784 3952 10836 4004
rect 22100 3952 22152 4004
rect 22192 3952 22244 4004
rect 23664 3995 23716 4004
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 9772 3884 9824 3936
rect 11336 3884 11388 3936
rect 16028 3884 16080 3936
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 18972 3927 19024 3936
rect 18972 3893 18981 3927
rect 18981 3893 19015 3927
rect 19015 3893 19024 3927
rect 18972 3884 19024 3893
rect 19064 3884 19116 3936
rect 20260 3884 20312 3936
rect 20352 3884 20404 3936
rect 23664 3961 23673 3995
rect 23673 3961 23707 3995
rect 23707 3961 23716 3995
rect 23664 3952 23716 3961
rect 29000 4088 29052 4140
rect 30288 4088 30340 4140
rect 29552 4020 29604 4072
rect 36084 4156 36136 4208
rect 31944 4088 31996 4140
rect 32128 4088 32180 4140
rect 33784 4088 33836 4140
rect 33048 4020 33100 4072
rect 35900 4020 35952 4072
rect 37832 4088 37884 4140
rect 40776 4156 40828 4208
rect 38384 4088 38436 4140
rect 38568 4131 38620 4140
rect 38568 4097 38577 4131
rect 38577 4097 38611 4131
rect 38611 4097 38620 4131
rect 38568 4088 38620 4097
rect 38752 4088 38804 4140
rect 41052 4088 41104 4140
rect 41236 4088 41288 4140
rect 43812 4233 43821 4267
rect 43821 4233 43855 4267
rect 43855 4233 43864 4267
rect 43812 4224 43864 4233
rect 45468 4224 45520 4276
rect 46388 4156 46440 4208
rect 25964 3884 26016 3936
rect 26424 3884 26476 3936
rect 26884 3884 26936 3936
rect 33784 3952 33836 4004
rect 35808 3952 35860 4004
rect 36636 3952 36688 4004
rect 38752 3952 38804 4004
rect 40868 3952 40920 4004
rect 29552 3884 29604 3936
rect 30196 3884 30248 3936
rect 32128 3884 32180 3936
rect 32496 3927 32548 3936
rect 32496 3893 32505 3927
rect 32505 3893 32539 3927
rect 32539 3893 32548 3927
rect 32496 3884 32548 3893
rect 32588 3884 32640 3936
rect 35348 3884 35400 3936
rect 36452 3884 36504 3936
rect 38844 3927 38896 3936
rect 38844 3893 38853 3927
rect 38853 3893 38887 3927
rect 38887 3893 38896 3927
rect 38844 3884 38896 3893
rect 40960 3884 41012 3936
rect 41328 3952 41380 4004
rect 41420 3952 41472 4004
rect 45468 4131 45520 4140
rect 45468 4097 45477 4131
rect 45477 4097 45511 4131
rect 45511 4097 45520 4131
rect 45468 4088 45520 4097
rect 45744 4131 45796 4140
rect 45744 4097 45753 4131
rect 45753 4097 45787 4131
rect 45787 4097 45796 4131
rect 45744 4088 45796 4097
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 48872 4224 48924 4276
rect 45836 4088 45888 4097
rect 41972 4020 42024 4072
rect 42432 4063 42484 4072
rect 42432 4029 42441 4063
rect 42441 4029 42475 4063
rect 42475 4029 42484 4063
rect 42432 4020 42484 4029
rect 47032 4156 47084 4208
rect 46848 4131 46900 4140
rect 46848 4097 46857 4131
rect 46857 4097 46891 4131
rect 46891 4097 46900 4131
rect 46848 4088 46900 4097
rect 47584 4131 47636 4140
rect 47584 4097 47593 4131
rect 47593 4097 47627 4131
rect 47627 4097 47636 4131
rect 47584 4088 47636 4097
rect 48688 4156 48740 4208
rect 48044 4088 48096 4140
rect 48780 4131 48832 4140
rect 48780 4097 48809 4131
rect 48809 4097 48832 4131
rect 49056 4131 49108 4140
rect 48780 4088 48832 4097
rect 49056 4097 49065 4131
rect 49065 4097 49099 4131
rect 49099 4097 49108 4131
rect 49056 4088 49108 4097
rect 49148 4131 49200 4140
rect 49148 4097 49157 4131
rect 49157 4097 49191 4131
rect 49191 4097 49200 4131
rect 49148 4088 49200 4097
rect 48044 3952 48096 4004
rect 49332 3995 49384 4004
rect 49332 3961 49341 3995
rect 49341 3961 49375 3995
rect 49375 3961 49384 3995
rect 49332 3952 49384 3961
rect 47032 3927 47084 3936
rect 47032 3893 47041 3927
rect 47041 3893 47075 3927
rect 47075 3893 47084 3927
rect 47032 3884 47084 3893
rect 47584 3884 47636 3936
rect 50160 3884 50212 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2964 3680 3016 3732
rect 5356 3680 5408 3732
rect 6644 3680 6696 3732
rect 7196 3723 7248 3732
rect 6736 3612 6788 3664
rect 6920 3612 6972 3664
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 7748 3680 7800 3732
rect 9128 3680 9180 3732
rect 10876 3680 10928 3732
rect 35900 3680 35952 3732
rect 36912 3723 36964 3732
rect 36912 3689 36921 3723
rect 36921 3689 36955 3723
rect 36955 3689 36964 3723
rect 36912 3680 36964 3689
rect 38384 3680 38436 3732
rect 39396 3680 39448 3732
rect 41420 3680 41472 3732
rect 42800 3723 42852 3732
rect 42800 3689 42809 3723
rect 42809 3689 42843 3723
rect 42843 3689 42852 3723
rect 42800 3680 42852 3689
rect 9312 3612 9364 3664
rect 9404 3612 9456 3664
rect 14924 3612 14976 3664
rect 16580 3612 16632 3664
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 9220 3544 9272 3596
rect 12992 3587 13044 3596
rect 204 3408 256 3460
rect 5080 3476 5132 3528
rect 5264 3476 5316 3528
rect 5540 3476 5592 3528
rect 6736 3476 6788 3528
rect 7472 3476 7524 3528
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 9496 3519 9548 3528
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9680 3519 9732 3528
rect 9496 3476 9548 3485
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 10600 3519 10652 3528
rect 9772 3476 9824 3485
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 13912 3544 13964 3596
rect 15476 3587 15528 3596
rect 3608 3340 3660 3392
rect 4620 3383 4672 3392
rect 4620 3349 4629 3383
rect 4629 3349 4663 3383
rect 4663 3349 4672 3383
rect 4620 3340 4672 3349
rect 5080 3340 5132 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 8668 3340 8720 3392
rect 10876 3408 10928 3460
rect 14004 3476 14056 3528
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 15752 3519 15804 3528
rect 15752 3485 15786 3519
rect 15786 3485 15804 3519
rect 15752 3476 15804 3485
rect 20168 3612 20220 3664
rect 21824 3612 21876 3664
rect 22100 3612 22152 3664
rect 22192 3612 22244 3664
rect 23020 3612 23072 3664
rect 23296 3655 23348 3664
rect 23296 3621 23305 3655
rect 23305 3621 23339 3655
rect 23339 3621 23348 3655
rect 23296 3612 23348 3621
rect 24492 3612 24544 3664
rect 20352 3544 20404 3596
rect 24400 3544 24452 3596
rect 18788 3476 18840 3528
rect 20260 3476 20312 3528
rect 20536 3476 20588 3528
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 22744 3519 22796 3528
rect 22744 3485 22754 3519
rect 22754 3485 22788 3519
rect 22788 3485 22796 3519
rect 23020 3519 23072 3528
rect 22744 3476 22796 3485
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 23480 3476 23532 3528
rect 24492 3476 24544 3528
rect 24860 3519 24912 3528
rect 24860 3485 24873 3519
rect 24873 3485 24907 3519
rect 24907 3485 24912 3519
rect 24860 3476 24912 3485
rect 13360 3408 13412 3460
rect 17132 3408 17184 3460
rect 10784 3340 10836 3392
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 15384 3340 15436 3392
rect 15476 3340 15528 3392
rect 17316 3340 17368 3392
rect 17684 3340 17736 3392
rect 18512 3383 18564 3392
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 19248 3383 19300 3392
rect 19248 3349 19257 3383
rect 19257 3349 19291 3383
rect 19291 3349 19300 3383
rect 19248 3340 19300 3349
rect 21088 3408 21140 3460
rect 22928 3451 22980 3460
rect 22928 3417 22937 3451
rect 22937 3417 22971 3451
rect 22971 3417 22980 3451
rect 22928 3408 22980 3417
rect 23020 3340 23072 3392
rect 25872 3612 25924 3664
rect 26976 3612 27028 3664
rect 31208 3544 31260 3596
rect 36446 3587 36498 3596
rect 25596 3476 25648 3528
rect 26424 3476 26476 3528
rect 31116 3476 31168 3528
rect 36446 3553 36455 3587
rect 36455 3553 36489 3587
rect 36489 3553 36498 3587
rect 36446 3544 36498 3553
rect 36728 3612 36780 3664
rect 43444 3612 43496 3664
rect 46388 3612 46440 3664
rect 47584 3680 47636 3732
rect 57152 3680 57204 3732
rect 47952 3612 48004 3664
rect 42156 3544 42208 3596
rect 47584 3544 47636 3596
rect 48504 3544 48556 3596
rect 31576 3476 31628 3528
rect 32128 3519 32180 3528
rect 32128 3485 32137 3519
rect 32137 3485 32171 3519
rect 32171 3485 32180 3519
rect 32128 3476 32180 3485
rect 25780 3408 25832 3460
rect 31208 3451 31260 3460
rect 31208 3417 31217 3451
rect 31217 3417 31251 3451
rect 31251 3417 31260 3451
rect 31208 3408 31260 3417
rect 25412 3383 25464 3392
rect 25412 3349 25421 3383
rect 25421 3349 25455 3383
rect 25455 3349 25464 3383
rect 25412 3340 25464 3349
rect 25964 3340 26016 3392
rect 31116 3340 31168 3392
rect 31576 3383 31628 3392
rect 31576 3349 31585 3383
rect 31585 3349 31619 3383
rect 31619 3349 31628 3383
rect 31576 3340 31628 3349
rect 34428 3408 34480 3460
rect 32312 3340 32364 3392
rect 34520 3340 34572 3392
rect 34796 3476 34848 3528
rect 35348 3476 35400 3528
rect 36084 3476 36136 3528
rect 35532 3408 35584 3460
rect 36636 3476 36688 3528
rect 37004 3476 37056 3528
rect 38200 3519 38252 3528
rect 38200 3485 38209 3519
rect 38209 3485 38243 3519
rect 38243 3485 38252 3519
rect 38200 3476 38252 3485
rect 38292 3476 38344 3528
rect 40132 3476 40184 3528
rect 40776 3476 40828 3528
rect 41236 3519 41288 3528
rect 41236 3485 41245 3519
rect 41245 3485 41279 3519
rect 41279 3485 41288 3519
rect 41236 3476 41288 3485
rect 41512 3519 41564 3528
rect 41512 3485 41521 3519
rect 41521 3485 41555 3519
rect 41555 3485 41564 3519
rect 41512 3476 41564 3485
rect 42248 3519 42300 3528
rect 39856 3408 39908 3460
rect 41328 3408 41380 3460
rect 42248 3485 42257 3519
rect 42257 3485 42291 3519
rect 42291 3485 42300 3519
rect 42248 3476 42300 3485
rect 42524 3519 42576 3528
rect 42524 3485 42529 3519
rect 42529 3485 42563 3519
rect 42563 3485 42576 3519
rect 42524 3476 42576 3485
rect 42708 3476 42760 3528
rect 42800 3476 42852 3528
rect 43812 3476 43864 3528
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 45928 3519 45980 3528
rect 45928 3485 45937 3519
rect 45937 3485 45971 3519
rect 45971 3485 45980 3519
rect 45928 3476 45980 3485
rect 46296 3519 46348 3528
rect 39580 3340 39632 3392
rect 39672 3340 39724 3392
rect 40868 3340 40920 3392
rect 46296 3485 46305 3519
rect 46305 3485 46339 3519
rect 46339 3485 46348 3519
rect 46296 3476 46348 3485
rect 46940 3519 46992 3528
rect 46940 3485 46949 3519
rect 46949 3485 46983 3519
rect 46983 3485 46992 3519
rect 46940 3476 46992 3485
rect 47124 3519 47176 3528
rect 47124 3485 47133 3519
rect 47133 3485 47167 3519
rect 47167 3485 47176 3519
rect 47124 3476 47176 3485
rect 47492 3476 47544 3528
rect 47860 3476 47912 3528
rect 48872 3476 48924 3528
rect 51172 3544 51224 3596
rect 41788 3383 41840 3392
rect 41788 3349 41797 3383
rect 41797 3349 41831 3383
rect 41831 3349 41840 3383
rect 41788 3340 41840 3349
rect 42708 3340 42760 3392
rect 46664 3408 46716 3460
rect 47216 3451 47268 3460
rect 47216 3417 47225 3451
rect 47225 3417 47259 3451
rect 47259 3417 47268 3451
rect 47216 3408 47268 3417
rect 48044 3408 48096 3460
rect 49608 3476 49660 3528
rect 58164 3476 58216 3528
rect 42984 3340 43036 3392
rect 45468 3340 45520 3392
rect 46480 3383 46532 3392
rect 46480 3349 46489 3383
rect 46489 3349 46523 3383
rect 46523 3349 46532 3383
rect 46480 3340 46532 3349
rect 46940 3340 46992 3392
rect 48320 3340 48372 3392
rect 48412 3340 48464 3392
rect 51540 3383 51592 3392
rect 51540 3349 51549 3383
rect 51549 3349 51583 3383
rect 51583 3349 51592 3383
rect 51540 3340 51592 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 3240 3000 3292 3052
rect 5172 3068 5224 3120
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6828 3068 6880 3120
rect 8300 3136 8352 3188
rect 8392 3136 8444 3188
rect 9404 3111 9456 3120
rect 1952 2932 2004 2984
rect 3332 2932 3384 2984
rect 3792 2932 3844 2984
rect 5448 2932 5500 2984
rect 664 2864 716 2916
rect 7564 3000 7616 3052
rect 8392 3000 8444 3052
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 9404 3077 9438 3111
rect 9438 3077 9456 3111
rect 9404 3068 9456 3077
rect 9588 3136 9640 3188
rect 15108 3136 15160 3188
rect 9956 3000 10008 3052
rect 10968 3000 11020 3052
rect 12992 3000 13044 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 2596 2796 2648 2848
rect 4712 2796 4764 2848
rect 7288 2864 7340 2916
rect 10140 2932 10192 2984
rect 19340 3136 19392 3188
rect 19984 3136 20036 3188
rect 20076 3136 20128 3188
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 22376 3136 22428 3188
rect 24860 3136 24912 3188
rect 17316 3068 17368 3120
rect 16028 3043 16080 3052
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 17500 3000 17552 3052
rect 18972 3068 19024 3120
rect 22008 3068 22060 3120
rect 23020 3111 23072 3120
rect 20260 3000 20312 3052
rect 21088 3000 21140 3052
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 22652 3043 22704 3052
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 23020 3077 23029 3111
rect 23029 3077 23063 3111
rect 23063 3077 23072 3111
rect 23020 3068 23072 3077
rect 25596 3136 25648 3188
rect 25688 3136 25740 3188
rect 27252 3136 27304 3188
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 23480 3000 23532 3052
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 24124 3000 24176 3052
rect 25412 3068 25464 3120
rect 31024 3136 31076 3188
rect 31208 3136 31260 3188
rect 31852 3136 31904 3188
rect 31392 3068 31444 3120
rect 33876 3068 33928 3120
rect 34704 3136 34756 3188
rect 39396 3136 39448 3188
rect 39856 3136 39908 3188
rect 41328 3179 41380 3188
rect 41328 3145 41337 3179
rect 41337 3145 41371 3179
rect 41371 3145 41380 3179
rect 41328 3136 41380 3145
rect 36912 3068 36964 3120
rect 22468 2932 22520 2984
rect 25964 3000 26016 3052
rect 27436 3000 27488 3052
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 30840 3000 30892 3052
rect 31116 3043 31168 3052
rect 31116 3009 31125 3043
rect 31125 3009 31159 3043
rect 31159 3009 31168 3043
rect 31116 3000 31168 3009
rect 32404 3043 32456 3052
rect 14832 2864 14884 2916
rect 30288 2932 30340 2984
rect 32404 3009 32413 3043
rect 32413 3009 32447 3043
rect 32447 3009 32456 3043
rect 32404 3000 32456 3009
rect 33416 3043 33468 3052
rect 33416 3009 33425 3043
rect 33425 3009 33459 3043
rect 33459 3009 33468 3043
rect 33416 3000 33468 3009
rect 31944 2932 31996 2984
rect 32312 2932 32364 2984
rect 34520 3000 34572 3052
rect 38844 3068 38896 3120
rect 41052 3111 41104 3120
rect 41052 3077 41061 3111
rect 41061 3077 41095 3111
rect 41095 3077 41104 3111
rect 42248 3136 42300 3188
rect 48688 3136 48740 3188
rect 41052 3068 41104 3077
rect 41788 3068 41840 3120
rect 47032 3068 47084 3120
rect 49608 3068 49660 3120
rect 38108 3000 38160 3052
rect 38292 3000 38344 3052
rect 35256 2975 35308 2984
rect 35256 2941 35265 2975
rect 35265 2941 35299 2975
rect 35299 2941 35308 2975
rect 35256 2932 35308 2941
rect 37924 2932 37976 2984
rect 39856 3000 39908 3052
rect 40776 3043 40828 3052
rect 40776 3009 40785 3043
rect 40785 3009 40819 3043
rect 40819 3009 40828 3043
rect 40776 3000 40828 3009
rect 40868 3000 40920 3052
rect 41144 3043 41196 3052
rect 41144 3009 41153 3043
rect 41153 3009 41187 3043
rect 41187 3009 41196 3043
rect 41144 3000 41196 3009
rect 43904 3000 43956 3052
rect 45652 3043 45704 3052
rect 45652 3009 45661 3043
rect 45661 3009 45695 3043
rect 45695 3009 45704 3043
rect 45652 3000 45704 3009
rect 45928 3043 45980 3052
rect 45928 3009 45962 3043
rect 45962 3009 45980 3043
rect 45928 3000 45980 3009
rect 47768 3000 47820 3052
rect 48596 3000 48648 3052
rect 50160 3000 50212 3052
rect 52184 3000 52236 3052
rect 55864 3043 55916 3052
rect 42432 2975 42484 2984
rect 5448 2796 5500 2848
rect 9772 2796 9824 2848
rect 12256 2796 12308 2848
rect 15108 2796 15160 2848
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 16764 2796 16816 2848
rect 17224 2796 17276 2848
rect 22652 2864 22704 2916
rect 21640 2796 21692 2848
rect 22928 2796 22980 2848
rect 23756 2796 23808 2848
rect 25136 2796 25188 2848
rect 25596 2796 25648 2848
rect 25872 2796 25924 2848
rect 30288 2796 30340 2848
rect 32312 2796 32364 2848
rect 37004 2864 37056 2916
rect 36728 2796 36780 2848
rect 38200 2796 38252 2848
rect 42432 2941 42441 2975
rect 42441 2941 42475 2975
rect 42475 2941 42484 2975
rect 42432 2932 42484 2941
rect 46756 2932 46808 2984
rect 41144 2864 41196 2916
rect 46940 2864 46992 2916
rect 42616 2796 42668 2848
rect 44088 2796 44140 2848
rect 45652 2796 45704 2848
rect 46388 2796 46440 2848
rect 46664 2796 46716 2848
rect 48780 2796 48832 2848
rect 51540 2932 51592 2984
rect 55864 3009 55873 3043
rect 55873 3009 55907 3043
rect 55907 3009 55916 3043
rect 55864 3000 55916 3009
rect 59636 3136 59688 3188
rect 57152 3111 57204 3120
rect 57152 3077 57161 3111
rect 57161 3077 57195 3111
rect 57195 3077 57204 3111
rect 57152 3068 57204 3077
rect 50160 2864 50212 2916
rect 51356 2796 51408 2848
rect 52828 2796 52880 2848
rect 54300 2796 54352 2848
rect 55772 2796 55824 2848
rect 58716 2796 58768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3700 2592 3752 2644
rect 4896 2592 4948 2644
rect 1124 2524 1176 2576
rect 5540 2524 5592 2576
rect 3332 2456 3384 2508
rect 6276 2456 6328 2508
rect 4620 2388 4672 2440
rect 8852 2456 8904 2508
rect 7104 2431 7156 2440
rect 1308 2320 1360 2372
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 11888 2592 11940 2644
rect 9404 2524 9456 2576
rect 12348 2524 12400 2576
rect 19340 2592 19392 2644
rect 22192 2592 22244 2644
rect 22468 2592 22520 2644
rect 22836 2592 22888 2644
rect 25596 2592 25648 2644
rect 28908 2592 28960 2644
rect 30104 2592 30156 2644
rect 34612 2592 34664 2644
rect 9772 2388 9824 2440
rect 12256 2431 12308 2440
rect 8760 2320 8812 2372
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 15292 2456 15344 2508
rect 15108 2431 15160 2440
rect 15108 2397 15117 2431
rect 15117 2397 15151 2431
rect 15151 2397 15160 2431
rect 15108 2388 15160 2397
rect 17132 2388 17184 2440
rect 17316 2388 17368 2440
rect 18512 2388 18564 2440
rect 22100 2524 22152 2576
rect 25044 2524 25096 2576
rect 20904 2456 20956 2508
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 3056 2252 3108 2304
rect 6000 2252 6052 2304
rect 6736 2252 6788 2304
rect 7932 2252 7984 2304
rect 8484 2252 8536 2304
rect 9220 2252 9272 2304
rect 11336 2252 11388 2304
rect 11888 2252 11940 2304
rect 14280 2252 14332 2304
rect 14832 2252 14884 2304
rect 15384 2252 15436 2304
rect 19064 2320 19116 2372
rect 22928 2388 22980 2440
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 24308 2320 24360 2372
rect 24860 2388 24912 2440
rect 26884 2388 26936 2440
rect 30840 2524 30892 2576
rect 32956 2524 33008 2576
rect 30288 2456 30340 2508
rect 31484 2456 31536 2508
rect 33324 2456 33376 2508
rect 35624 2592 35676 2644
rect 45928 2592 45980 2644
rect 37004 2524 37056 2576
rect 49056 2524 49108 2576
rect 41328 2456 41380 2508
rect 51264 2499 51316 2508
rect 51264 2465 51273 2499
rect 51273 2465 51307 2499
rect 51307 2465 51316 2499
rect 51264 2456 51316 2465
rect 52644 2456 52696 2508
rect 28264 2388 28316 2440
rect 28908 2388 28960 2440
rect 29552 2431 29604 2440
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 30380 2388 30432 2440
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31852 2388 31904 2440
rect 34428 2388 34480 2440
rect 34704 2320 34756 2372
rect 36268 2388 36320 2440
rect 37556 2431 37608 2440
rect 37556 2397 37565 2431
rect 37565 2397 37599 2431
rect 37599 2397 37608 2431
rect 37556 2388 37608 2397
rect 37096 2320 37148 2372
rect 45376 2388 45428 2440
rect 45652 2431 45704 2440
rect 45652 2397 45661 2431
rect 45661 2397 45695 2431
rect 45695 2397 45704 2431
rect 45652 2388 45704 2397
rect 45836 2431 45888 2440
rect 45836 2397 45845 2431
rect 45845 2397 45879 2431
rect 45879 2397 45888 2431
rect 45836 2388 45888 2397
rect 47952 2388 48004 2440
rect 49424 2388 49476 2440
rect 50896 2388 50948 2440
rect 52368 2388 52420 2440
rect 53840 2388 53892 2440
rect 55220 2388 55272 2440
rect 56692 2388 56744 2440
rect 37740 2320 37792 2372
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 42064 2320 42116 2372
rect 43536 2320 43588 2372
rect 45744 2363 45796 2372
rect 45744 2329 45753 2363
rect 45753 2329 45787 2363
rect 45787 2329 45796 2363
rect 45744 2320 45796 2329
rect 19156 2252 19208 2304
rect 19984 2252 20036 2304
rect 20536 2252 20588 2304
rect 24032 2252 24084 2304
rect 24676 2252 24728 2304
rect 26516 2252 26568 2304
rect 27988 2252 28040 2304
rect 29460 2252 29512 2304
rect 30840 2252 30892 2304
rect 33784 2252 33836 2304
rect 35256 2252 35308 2304
rect 36544 2252 36596 2304
rect 37832 2252 37884 2304
rect 38752 2295 38804 2304
rect 38752 2261 38761 2295
rect 38761 2261 38795 2295
rect 38795 2261 38804 2295
rect 38752 2252 38804 2261
rect 45008 2252 45060 2304
rect 46756 2320 46808 2372
rect 48228 2320 48280 2372
rect 53012 2363 53064 2372
rect 53012 2329 53021 2363
rect 53021 2329 53055 2363
rect 53055 2329 53064 2363
rect 53012 2320 53064 2329
rect 54208 2363 54260 2372
rect 54208 2329 54217 2363
rect 54217 2329 54251 2363
rect 54251 2329 54260 2363
rect 54208 2320 54260 2329
rect 55588 2363 55640 2372
rect 55588 2329 55597 2363
rect 55597 2329 55631 2363
rect 55631 2329 55640 2363
rect 55588 2320 55640 2329
rect 57060 2363 57112 2372
rect 57060 2329 57069 2363
rect 57069 2329 57103 2363
rect 57103 2329 57112 2363
rect 57060 2320 57112 2329
rect 48136 2295 48188 2304
rect 48136 2261 48145 2295
rect 48145 2261 48179 2295
rect 48179 2261 48188 2295
rect 48136 2252 48188 2261
rect 48872 2295 48924 2304
rect 48872 2261 48881 2295
rect 48881 2261 48915 2295
rect 48915 2261 48924 2295
rect 48872 2252 48924 2261
rect 57244 2252 57296 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 6368 2048 6420 2100
rect 23204 2048 23256 2100
rect 26884 2048 26936 2100
rect 32036 2048 32088 2100
rect 37188 2048 37240 2100
rect 41328 2048 41380 2100
rect 12992 1980 13044 2032
rect 22008 1980 22060 2032
rect 31668 1980 31720 2032
rect 37556 1980 37608 2032
rect 37832 1980 37884 2032
rect 48136 1980 48188 2032
rect 16304 1912 16356 1964
rect 57060 1912 57112 1964
rect 20444 1844 20496 1896
rect 45744 1844 45796 1896
rect 16396 1776 16448 1828
rect 55588 1776 55640 1828
rect 12716 1708 12768 1760
rect 54208 1708 54260 1760
rect 10232 1640 10284 1692
rect 48228 1640 48280 1692
rect 10692 1572 10744 1624
rect 53012 1572 53064 1624
rect 37648 1504 37700 1556
rect 48872 1504 48924 1556
rect 7104 1436 7156 1488
rect 22744 1436 22796 1488
rect 33508 1436 33560 1488
rect 38752 1436 38804 1488
rect 3332 1028 3384 1080
rect 8576 1028 8628 1080
<< metal2 >>
rect 2962 41712 3018 41721
rect 2962 41647 3018 41656
rect 2778 40080 2834 40089
rect 2778 40015 2834 40024
rect 2792 39642 2820 40015
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 1768 39432 1820 39438
rect 1768 39374 1820 39380
rect 2320 39432 2372 39438
rect 2320 39374 2372 39380
rect 2872 39432 2924 39438
rect 2872 39374 2924 39380
rect 1584 39296 1636 39302
rect 1582 39264 1584 39273
rect 1636 39264 1638 39273
rect 1582 39199 1638 39208
rect 1584 38752 1636 38758
rect 1584 38694 1636 38700
rect 1596 38457 1624 38694
rect 1582 38448 1638 38457
rect 1582 38383 1638 38392
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 1584 37664 1636 37670
rect 1582 37632 1584 37641
rect 1636 37632 1638 37641
rect 1582 37567 1638 37576
rect 1582 36680 1638 36689
rect 1582 36615 1584 36624
rect 1636 36615 1638 36624
rect 1584 36586 1636 36592
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35873 1624 35974
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 1582 35048 1638 35057
rect 1582 34983 1638 34992
rect 1596 34746 1624 34983
rect 1584 34740 1636 34746
rect 1584 34682 1636 34688
rect 1584 33856 1636 33862
rect 1582 33824 1584 33833
rect 1636 33824 1638 33833
rect 1582 33759 1638 33768
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 33425 1440 33458
rect 1398 33416 1454 33425
rect 1398 33351 1454 33360
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1596 32473 1624 32710
rect 1582 32464 1638 32473
rect 1400 32428 1452 32434
rect 1582 32399 1638 32408
rect 1400 32370 1452 32376
rect 1412 32065 1440 32370
rect 1398 32056 1454 32065
rect 1398 31991 1454 32000
rect 1584 31680 1636 31686
rect 1584 31622 1636 31628
rect 1596 31249 1624 31622
rect 1582 31240 1638 31249
rect 1582 31175 1638 31184
rect 1688 31090 1716 37810
rect 1780 35170 1808 39374
rect 2044 36168 2096 36174
rect 2044 36110 2096 36116
rect 2056 35894 2084 36110
rect 2332 35894 2360 39374
rect 2884 35894 2912 39374
rect 2976 38554 3004 41647
rect 3698 41200 3754 42000
rect 11150 41200 11206 42000
rect 18694 41200 18750 42000
rect 26146 41200 26202 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48686 41200 48742 42000
rect 56138 41200 56194 42000
rect 3054 40896 3110 40905
rect 3054 40831 3110 40840
rect 3068 39642 3096 40831
rect 3712 39642 3740 41200
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 3056 39636 3108 39642
rect 3056 39578 3108 39584
rect 3700 39636 3752 39642
rect 3700 39578 3752 39584
rect 18708 39506 18736 41200
rect 26160 39658 26188 41200
rect 26160 39642 26280 39658
rect 26160 39636 26292 39642
rect 26160 39630 26240 39636
rect 26240 39578 26292 39584
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 33704 39438 33732 41200
rect 41156 39930 41184 41200
rect 41156 39902 41460 39930
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 41432 39642 41460 39902
rect 48700 39642 48728 41200
rect 56152 39642 56180 41200
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 48688 39636 48740 39642
rect 48688 39578 48740 39584
rect 56140 39636 56192 39642
rect 56140 39578 56192 39584
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 32128 39432 32180 39438
rect 32128 39374 32180 39380
rect 33692 39432 33744 39438
rect 33692 39374 33744 39380
rect 54760 39432 54812 39438
rect 54760 39374 54812 39380
rect 2964 38548 3016 38554
rect 2964 38490 3016 38496
rect 2056 35866 2176 35894
rect 2332 35866 2636 35894
rect 2884 35866 3004 35894
rect 1780 35142 2084 35170
rect 1860 35012 1912 35018
rect 1860 34954 1912 34960
rect 1872 34649 1900 34954
rect 1952 34944 2004 34950
rect 1952 34886 2004 34892
rect 1858 34640 1914 34649
rect 1858 34575 1914 34584
rect 1768 31340 1820 31346
rect 1768 31282 1820 31288
rect 1504 31062 1716 31090
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1412 29209 1440 30194
rect 1398 29200 1454 29209
rect 1398 29135 1454 29144
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27130 1440 28018
rect 1400 27124 1452 27130
rect 1400 27066 1452 27072
rect 1400 26920 1452 26926
rect 1400 26862 1452 26868
rect 1412 24750 1440 26862
rect 1504 24750 1532 31062
rect 1780 30841 1808 31282
rect 1766 30832 1822 30841
rect 1766 30767 1822 30776
rect 1584 30592 1636 30598
rect 1584 30534 1636 30540
rect 1596 30025 1624 30534
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1676 29640 1728 29646
rect 1674 29608 1676 29617
rect 1728 29608 1730 29617
rect 1674 29543 1730 29552
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28801 1624 28970
rect 1582 28792 1638 28801
rect 1582 28727 1638 28736
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 27441 1624 27814
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1584 26240 1636 26246
rect 1582 26208 1584 26217
rect 1636 26208 1638 26217
rect 1582 26143 1638 26152
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24993 1624 25094
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1688 24886 1716 29242
rect 1872 29102 1900 30126
rect 1860 29096 1912 29102
rect 1860 29038 1912 29044
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 1768 28416 1820 28422
rect 1872 28393 1900 28426
rect 1768 28358 1820 28364
rect 1858 28384 1914 28393
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1490 24576 1546 24585
rect 1412 24274 1440 24550
rect 1490 24511 1546 24520
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1504 24206 1532 24511
rect 1492 24200 1544 24206
rect 1596 24177 1624 24754
rect 1676 24744 1728 24750
rect 1676 24686 1728 24692
rect 1492 24142 1544 24148
rect 1582 24168 1638 24177
rect 1688 24138 1716 24686
rect 1780 24154 1808 28358
rect 1858 28319 1914 28328
rect 1860 27396 1912 27402
rect 1860 27338 1912 27344
rect 1872 27033 1900 27338
rect 1858 27024 1914 27033
rect 1858 26959 1914 26968
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1872 25809 1900 25842
rect 1858 25800 1914 25809
rect 1858 25735 1914 25744
rect 1582 24103 1638 24112
rect 1676 24132 1728 24138
rect 1780 24126 1900 24154
rect 1676 24074 1728 24080
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1596 23769 1624 23802
rect 1582 23760 1638 23769
rect 1582 23695 1638 23704
rect 1780 23526 1808 24006
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1398 23216 1454 23225
rect 1398 23151 1400 23160
rect 1452 23151 1454 23160
rect 1400 23122 1452 23128
rect 1676 23112 1728 23118
rect 1676 23054 1728 23060
rect 1688 22710 1716 23054
rect 1676 22704 1728 22710
rect 1676 22646 1728 22652
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22234 1440 22578
rect 1492 22500 1544 22506
rect 1492 22442 1544 22448
rect 1400 22228 1452 22234
rect 1400 22170 1452 22176
rect 1504 21010 1532 22442
rect 1584 22432 1636 22438
rect 1582 22400 1584 22409
rect 1636 22400 1638 22409
rect 1582 22335 1638 22344
rect 1872 22250 1900 24126
rect 1780 22222 1900 22250
rect 1780 21706 1808 22222
rect 1860 22024 1912 22030
rect 1858 21992 1860 22001
rect 1912 21992 1914 22001
rect 1858 21927 1914 21936
rect 1688 21678 1808 21706
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1504 19922 1532 20946
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19961 1624 20198
rect 1582 19952 1638 19961
rect 1492 19916 1544 19922
rect 1582 19887 1638 19896
rect 1492 19858 1544 19864
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 17785 1440 19314
rect 1504 18766 1532 19858
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16153 1440 16934
rect 1504 16590 1532 18702
rect 1582 18592 1638 18601
rect 1582 18527 1638 18536
rect 1596 18426 1624 18527
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1688 17066 1716 21678
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 18630 1808 21490
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1872 19553 1900 19722
rect 1858 19544 1914 19553
rect 1858 19479 1914 19488
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1858 18184 1914 18193
rect 1858 18119 1914 18128
rect 1872 17678 1900 18119
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1964 17270 1992 34886
rect 2056 24070 2084 35142
rect 2148 29306 2176 35866
rect 2320 34604 2372 34610
rect 2320 34546 2372 34552
rect 2332 34241 2360 34546
rect 2318 34232 2374 34241
rect 2318 34167 2374 34176
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2136 29300 2188 29306
rect 2136 29242 2188 29248
rect 2136 29096 2188 29102
rect 2136 29038 2188 29044
rect 2148 28014 2176 29038
rect 2136 28008 2188 28014
rect 2136 27950 2188 27956
rect 2148 26790 2176 27950
rect 2136 26784 2188 26790
rect 2136 26726 2188 26732
rect 2136 25696 2188 25702
rect 2136 25638 2188 25644
rect 2148 25498 2176 25638
rect 2136 25492 2188 25498
rect 2136 25434 2188 25440
rect 2240 25378 2268 33390
rect 2320 31816 2372 31822
rect 2320 31758 2372 31764
rect 2332 31657 2360 31758
rect 2318 31648 2374 31657
rect 2318 31583 2374 31592
rect 2504 31272 2556 31278
rect 2504 31214 2556 31220
rect 2412 30728 2464 30734
rect 2412 30670 2464 30676
rect 2320 30592 2372 30598
rect 2320 30534 2372 30540
rect 2332 30258 2360 30534
rect 2320 30252 2372 30258
rect 2320 30194 2372 30200
rect 2318 30152 2374 30161
rect 2318 30087 2374 30096
rect 2332 27606 2360 30087
rect 2424 29850 2452 30670
rect 2412 29844 2464 29850
rect 2412 29786 2464 29792
rect 2320 27600 2372 27606
rect 2320 27542 2372 27548
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2332 26586 2360 27406
rect 2320 26580 2372 26586
rect 2320 26522 2372 26528
rect 2148 25350 2268 25378
rect 2516 25378 2544 31214
rect 2608 30161 2636 35866
rect 2780 33516 2832 33522
rect 2780 33458 2832 33464
rect 2792 33017 2820 33458
rect 2778 33008 2834 33017
rect 2778 32943 2834 32952
rect 2688 30592 2740 30598
rect 2688 30534 2740 30540
rect 2594 30152 2650 30161
rect 2594 30087 2650 30096
rect 2596 29776 2648 29782
rect 2596 29718 2648 29724
rect 2608 28626 2636 29718
rect 2700 29714 2728 30534
rect 2688 29708 2740 29714
rect 2688 29650 2740 29656
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2596 28620 2648 28626
rect 2596 28562 2648 28568
rect 2608 26518 2636 28562
rect 2700 28218 2728 29106
rect 2780 29028 2832 29034
rect 2780 28970 2832 28976
rect 2688 28212 2740 28218
rect 2688 28154 2740 28160
rect 2792 28150 2820 28970
rect 2884 28762 2912 29106
rect 2872 28756 2924 28762
rect 2872 28698 2924 28704
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2688 27328 2740 27334
rect 2688 27270 2740 27276
rect 2780 27328 2832 27334
rect 2780 27270 2832 27276
rect 2700 27062 2728 27270
rect 2688 27056 2740 27062
rect 2688 26998 2740 27004
rect 2596 26512 2648 26518
rect 2596 26454 2648 26460
rect 2608 26042 2636 26454
rect 2792 26450 2820 27270
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2872 25900 2924 25906
rect 2872 25842 2924 25848
rect 2884 25401 2912 25842
rect 2976 25702 3004 35866
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 3068 30433 3096 30670
rect 3054 30424 3110 30433
rect 3054 30359 3110 30368
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 3424 30048 3476 30054
rect 3424 29990 3476 29996
rect 3068 28490 3096 29990
rect 3436 29578 3464 29990
rect 3424 29572 3476 29578
rect 3424 29514 3476 29520
rect 3332 29504 3384 29510
rect 3332 29446 3384 29452
rect 3056 28484 3108 28490
rect 3056 28426 3108 28432
rect 3344 27826 3372 29446
rect 3884 28416 3936 28422
rect 3884 28358 3936 28364
rect 3896 27946 3924 28358
rect 3884 27940 3936 27946
rect 3884 27882 3936 27888
rect 3974 27840 4030 27849
rect 3344 27798 3464 27826
rect 3332 26852 3384 26858
rect 3332 26794 3384 26800
rect 3344 26314 3372 26794
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 2964 25696 3016 25702
rect 2964 25638 3016 25644
rect 2870 25392 2926 25401
rect 2516 25350 2636 25378
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 21554 2084 23462
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2148 21434 2176 25350
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2240 23730 2268 24754
rect 2332 23866 2360 25230
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 2424 24818 2452 25094
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2516 24410 2544 25230
rect 2504 24404 2556 24410
rect 2504 24346 2556 24352
rect 2412 24336 2464 24342
rect 2608 24290 2636 25350
rect 2870 25327 2926 25336
rect 2412 24278 2464 24284
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2228 23724 2280 23730
rect 2280 23684 2360 23712
rect 2228 23666 2280 23672
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22778 2268 23054
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2332 22506 2360 23684
rect 2424 22574 2452 24278
rect 2516 24262 2636 24290
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 2320 22500 2372 22506
rect 2320 22442 2372 22448
rect 2320 21956 2372 21962
rect 2320 21898 2372 21904
rect 2056 21406 2176 21434
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 2056 16794 2084 21406
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2240 20942 2268 21286
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2136 19780 2188 19786
rect 2136 19722 2188 19728
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 1492 16584 1544 16590
rect 1492 16526 1544 16532
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1596 15745 1624 16050
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1582 15736 1638 15745
rect 1582 15671 1638 15680
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 14929 1624 15302
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1398 14512 1454 14521
rect 1398 14447 1400 14456
rect 1452 14447 1454 14456
rect 1400 14418 1452 14424
rect 1872 13802 1900 15846
rect 1964 15162 1992 16526
rect 2148 15706 2176 19722
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2240 19145 2268 19314
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2332 16182 2360 21898
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2424 20602 2452 21490
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 2516 19938 2544 24262
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2608 23066 2636 23734
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2700 23322 2728 23666
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2608 23038 2820 23066
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2700 22778 2728 22918
rect 2792 22778 2820 23038
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2700 22166 2728 22510
rect 2688 22160 2740 22166
rect 2688 22102 2740 22108
rect 2700 20398 2728 22102
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2884 21593 2912 21966
rect 2870 21584 2926 21593
rect 2870 21519 2926 21528
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2884 21010 2912 21286
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 2964 20800 3016 20806
rect 3068 20777 3096 21490
rect 2964 20742 3016 20748
rect 3054 20768 3110 20777
rect 2976 20602 3004 20742
rect 3054 20703 3110 20712
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2778 20360 2834 20369
rect 2608 20058 2636 20334
rect 2778 20295 2834 20304
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2516 19910 2636 19938
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2424 16250 2452 17138
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 16590 2544 16934
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2608 15094 2636 19910
rect 2792 19854 2820 20295
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 3344 19378 3372 20402
rect 3436 20058 3464 27798
rect 3974 27775 4030 27784
rect 3988 27470 4016 27775
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3988 26625 4016 26930
rect 3974 26616 4030 26625
rect 3974 26551 4030 26560
rect 4080 26234 4108 39374
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 32140 39098 32168 39374
rect 43444 39296 43496 39302
rect 43444 39238 43496 39244
rect 32128 39092 32180 39098
rect 32128 39034 32180 39040
rect 13268 38956 13320 38962
rect 13268 38898 13320 38904
rect 32496 38956 32548 38962
rect 32496 38898 32548 38904
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 12072 36780 12124 36786
rect 12072 36722 12124 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 6184 34536 6236 34542
rect 6184 34478 6236 34484
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4988 32020 5040 32026
rect 4988 31962 5040 31968
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4724 30326 4752 30534
rect 4712 30320 4764 30326
rect 4712 30262 4764 30268
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4908 29850 4936 30670
rect 4896 29844 4948 29850
rect 4896 29786 4948 29792
rect 5000 29714 5028 31962
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 5816 30048 5868 30054
rect 5816 29990 5868 29996
rect 5092 29850 5120 29990
rect 5080 29844 5132 29850
rect 5080 29786 5132 29792
rect 4988 29708 5040 29714
rect 4988 29650 5040 29656
rect 5828 29646 5856 29990
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5816 29164 5868 29170
rect 5816 29106 5868 29112
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 5828 28762 5856 29106
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5724 27464 5776 27470
rect 5724 27406 5776 27412
rect 5828 27418 5856 27542
rect 5368 27130 5396 27406
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 3896 26206 4108 26234
rect 3516 24676 3568 24682
rect 3516 24618 3568 24624
rect 3528 24206 3556 24618
rect 3516 24200 3568 24206
rect 3516 24142 3568 24148
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3528 23050 3556 23462
rect 3516 23044 3568 23050
rect 3516 22986 3568 22992
rect 3528 22642 3556 22986
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3896 22094 3924 26206
rect 4540 26042 4568 26318
rect 5000 26042 5028 26726
rect 5736 26586 5764 27406
rect 5828 27390 6040 27418
rect 6196 27402 6224 34478
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6380 29306 6408 29514
rect 6368 29300 6420 29306
rect 6368 29242 6420 29248
rect 6380 28558 6408 29242
rect 6368 28552 6420 28558
rect 6368 28494 6420 28500
rect 5908 26852 5960 26858
rect 5908 26794 5960 26800
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 5724 25968 5776 25974
rect 5724 25910 5776 25916
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4632 25226 4660 25842
rect 5448 25764 5500 25770
rect 5448 25706 5500 25712
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4632 24138 4660 25162
rect 5460 24954 5488 25706
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5172 24744 5224 24750
rect 5172 24686 5224 24692
rect 5184 24274 5212 24686
rect 5644 24614 5672 25230
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3988 22817 4016 23054
rect 3974 22808 4030 22817
rect 3974 22743 4030 22752
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 3804 22066 3924 22094
rect 3804 21434 3832 22066
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3896 21554 3924 21830
rect 3988 21690 4016 22578
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3804 21406 4108 21434
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3620 19854 3648 20198
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18358 2728 19110
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3160 18426 3188 18906
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 2688 18352 2740 18358
rect 2688 18294 2740 18300
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2700 17105 2728 17614
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17377 2912 17478
rect 2870 17368 2926 17377
rect 2870 17303 2926 17312
rect 2686 17096 2742 17105
rect 2686 17031 2742 17040
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2792 16250 2820 16390
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 3068 16046 3096 18158
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3344 17678 3372 18022
rect 3804 17814 3832 18634
rect 3896 18426 3924 19246
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3896 18222 3924 18362
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3344 16969 3372 17138
rect 3330 16960 3386 16969
rect 3330 16895 3386 16904
rect 3976 16584 4028 16590
rect 3974 16552 3976 16561
rect 4028 16552 4030 16561
rect 3974 16487 4030 16496
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16114 3832 16390
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2700 14618 2728 14962
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2884 14414 2912 15574
rect 3068 15570 3096 15982
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2318 13968 2374 13977
rect 2318 13903 2320 13912
rect 2372 13903 2374 13912
rect 2320 13874 2372 13880
rect 3068 13870 3096 15506
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3528 14822 3556 15438
rect 3988 15337 4016 15438
rect 3974 15328 4030 15337
rect 3974 15263 4030 15272
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 3056 13728 3108 13734
rect 3056 13670 3108 13676
rect 1596 13569 1624 13670
rect 1582 13560 1638 13569
rect 1582 13495 1638 13504
rect 3068 13326 3096 13670
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 1872 13161 1900 13194
rect 1858 13152 1914 13161
rect 1858 13087 1914 13096
rect 1398 12744 1454 12753
rect 1398 12679 1454 12688
rect 1412 12238 1440 12679
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1596 11529 1624 11698
rect 1582 11520 1638 11529
rect 1582 11455 1638 11464
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1596 11121 1624 11222
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 2056 10674 2084 11698
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1596 10305 1624 10610
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1766 8936 1822 8945
rect 1412 8129 1440 8910
rect 1766 8871 1822 8880
rect 1780 8566 1808 8871
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 2056 8430 2084 10610
rect 2240 8498 2268 13194
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 2700 12442 2728 12786
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10674 2360 10950
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2424 10266 2452 11086
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1952 7880 2004 7886
rect 2056 7868 2084 8366
rect 2004 7840 2084 7868
rect 1952 7822 2004 7828
rect 1582 7712 1638 7721
rect 1582 7647 1638 7656
rect 1596 7546 1624 7647
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 2056 6934 2084 7840
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2044 6928 2096 6934
rect 2332 6905 2360 7346
rect 2044 6870 2096 6876
rect 2318 6896 2374 6905
rect 2318 6831 2374 6840
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6497 1440 6734
rect 1398 6488 1454 6497
rect 1398 6423 1454 6432
rect 1584 6112 1636 6118
rect 1582 6080 1584 6089
rect 1636 6080 1638 6089
rect 1582 6015 1638 6024
rect 2516 5778 2544 11494
rect 2608 10198 2636 12242
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2700 11898 2728 12038
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2884 11762 2912 12582
rect 3344 11937 3372 12786
rect 3330 11928 3386 11937
rect 3330 11863 3386 11872
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10713 3096 11086
rect 3528 10742 3556 14758
rect 3804 13394 3832 14962
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3804 11830 3832 13330
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3516 10736 3568 10742
rect 3054 10704 3110 10713
rect 3516 10678 3568 10684
rect 3054 10639 3110 10648
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2608 6254 2636 10134
rect 3436 10062 3464 10406
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9178 2728 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8537 2912 8910
rect 2870 8528 2926 8537
rect 2870 8463 2926 8472
rect 3252 8090 3280 9522
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 7313 3004 7346
rect 2962 7304 3018 7313
rect 2962 7239 3018 7248
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6458 2820 6734
rect 3252 6458 3280 7210
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 5778 2636 6190
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 1858 5672 1914 5681
rect 1858 5607 1914 5616
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1688 4622 1716 5306
rect 1872 5302 1900 5607
rect 1860 5296 1912 5302
rect 1860 5238 1912 5244
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 204 3460 256 3466
rect 204 3402 256 3408
rect 216 800 244 3402
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1124 2576 1176 2582
rect 1124 2518 1176 2524
rect 1136 800 1164 2518
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1320 649 1348 2314
rect 1596 800 1624 4422
rect 2792 4146 2820 5034
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4321 2912 4966
rect 2976 4729 3004 6258
rect 3620 5778 3648 10474
rect 3804 10130 3832 11766
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8566 3832 8774
rect 3988 8566 4016 12718
rect 4080 12374 4108 21406
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4632 18290 4660 24074
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5092 22438 5120 23666
rect 5736 23186 5764 25910
rect 5816 24676 5868 24682
rect 5816 24618 5868 24624
rect 5828 23662 5856 24618
rect 5816 23656 5868 23662
rect 5816 23598 5868 23604
rect 5828 23322 5856 23598
rect 5920 23322 5948 26794
rect 6012 26518 6040 27390
rect 6184 27396 6236 27402
rect 6184 27338 6236 27344
rect 6564 27130 6592 34682
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 6644 33312 6696 33318
rect 6644 33254 6696 33260
rect 6656 28626 6684 33254
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6748 28422 6776 29582
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6748 27946 6776 28358
rect 6736 27940 6788 27946
rect 6736 27882 6788 27888
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6656 26994 6684 27270
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6196 26586 6224 26726
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6000 26512 6052 26518
rect 6000 26454 6052 26460
rect 6196 24750 6224 26522
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 6380 25974 6408 26182
rect 6368 25968 6420 25974
rect 6368 25910 6420 25916
rect 6276 25152 6328 25158
rect 6276 25094 6328 25100
rect 6288 24818 6316 25094
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6184 24744 6236 24750
rect 6184 24686 6236 24692
rect 6196 24410 6224 24686
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6380 23798 6408 24550
rect 6368 23792 6420 23798
rect 6368 23734 6420 23740
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5920 23050 5948 23258
rect 6380 23118 6408 23462
rect 6656 23186 6684 26930
rect 6840 26926 6868 28562
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 25158 6868 26862
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 5908 23044 5960 23050
rect 5908 22986 5960 22992
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5092 22030 5120 22374
rect 6656 22030 6684 23122
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6932 21350 6960 23734
rect 7116 22642 7144 29446
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7024 21978 7052 22374
rect 7116 22098 7144 22578
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7024 21962 7144 21978
rect 7024 21956 7156 21962
rect 7024 21950 7104 21956
rect 7104 21898 7156 21904
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 7024 20942 7052 21830
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7116 21486 7144 21626
rect 7208 21554 7236 23666
rect 7300 21690 7328 28358
rect 9508 27130 9536 33934
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9048 26586 9076 26930
rect 9036 26580 9088 26586
rect 9036 26522 9088 26528
rect 9508 26382 9536 27066
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9496 26376 9548 26382
rect 9496 26318 9548 26324
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 8864 24410 8892 25230
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 8864 23662 8892 24346
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7392 22642 7420 22918
rect 7484 22642 7512 23462
rect 7656 23248 7708 23254
rect 7656 23190 7708 23196
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6840 19922 6868 20402
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6932 19786 6960 20742
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19446 5212 19654
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 6932 19378 6960 19722
rect 7024 19718 7052 20402
rect 7116 19854 7144 21422
rect 7300 21350 7328 21490
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7116 19378 7144 19790
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 6932 18834 6960 19314
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4264 15026 4292 15098
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4632 12238 4660 18226
rect 6184 18148 6236 18154
rect 6184 18090 6236 18096
rect 6196 17882 6224 18090
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4816 16046 4844 17614
rect 6196 17542 6224 17818
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15162 4844 15982
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4080 8838 4108 11154
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4908 10062 4936 16458
rect 6656 16250 6684 17070
rect 6748 16454 6776 17546
rect 6840 17338 6868 18566
rect 6932 18290 6960 18566
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6288 15706 6316 16050
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6656 15502 6684 16186
rect 6748 15502 6776 16390
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5644 15162 5672 15370
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5092 14618 5120 14962
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5184 13462 5212 13874
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5368 11626 5396 14350
rect 5644 14278 5672 15098
rect 6748 14414 6776 15438
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 5920 12442 5948 12854
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 4080 8362 4108 8774
rect 4264 8498 4292 8910
rect 4356 8634 4384 9046
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4632 7886 4660 8434
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3792 6928 3844 6934
rect 5460 6914 5488 12106
rect 6104 10266 6132 13942
rect 7024 13870 7052 14894
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6736 12096 6788 12102
rect 7024 12084 7052 13806
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 12238 7144 13194
rect 7208 12850 7236 13262
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12238 7236 12786
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7024 12056 7236 12084
rect 6736 12038 6788 12044
rect 6748 11830 6776 12038
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6184 11144 6236 11150
rect 6288 11132 6316 11698
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6236 11104 6316 11132
rect 6184 11086 6236 11092
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6104 9722 6132 10202
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 3792 6870 3844 6876
rect 5368 6886 5488 6914
rect 3804 6798 3832 6870
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 2976 4162 3004 4422
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2884 4134 3004 4162
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1858 3904 1914 3913
rect 1858 3839 1914 3848
rect 1872 3534 1900 3839
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 1873 1900 2994
rect 1964 2990 1992 4014
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1858 1864 1914 1873
rect 1858 1799 1914 1808
rect 2148 800 2176 3878
rect 2688 3528 2740 3534
rect 2686 3496 2688 3505
rect 2740 3496 2742 3505
rect 2686 3431 2742 3440
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 800 2636 2790
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 2884 241 2912 4134
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2976 3738 3004 4014
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 800 3096 2246
rect 3160 1465 3188 5646
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3344 4282 3372 5510
rect 3620 5234 3648 5510
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3804 4622 3832 6734
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6322 5212 6598
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5234 4292 5578
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4622 3924 4966
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3712 4146 3740 4490
rect 3804 4185 3832 4558
rect 3884 4208 3936 4214
rect 3790 4176 3846 4185
rect 3700 4140 3752 4146
rect 3884 4150 3936 4156
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 3790 4111 3846 4120
rect 3700 4082 3752 4088
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 3058 3280 3946
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3344 2514 3372 2926
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3146 1456 3202 1465
rect 3146 1391 3202 1400
rect 3332 1080 3384 1086
rect 3330 1048 3332 1057
rect 3384 1048 3386 1057
rect 3330 983 3386 992
rect 3620 800 3648 3334
rect 3804 2990 3832 4111
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3698 2680 3754 2689
rect 3698 2615 3700 2624
rect 3752 2615 3754 2624
rect 3700 2586 3752 2592
rect 3896 2281 3924 4150
rect 4172 4026 4200 4150
rect 4080 3998 4200 4026
rect 4080 3097 4108 3998
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4066 3088 4122 3097
rect 4066 3023 4122 3032
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4632 2446 4660 3334
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 3882 2272 3938 2281
rect 3882 2207 3938 2216
rect 4724 1442 4752 2790
rect 4908 2650 4936 5170
rect 5000 4214 5028 5170
rect 5184 4758 5212 5510
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 5184 4486 5212 4694
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 5080 4208 5132 4214
rect 5132 4156 5212 4162
rect 5080 4150 5212 4156
rect 5092 4134 5212 4150
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3534 5120 3946
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4540 1414 4752 1442
rect 4540 800 4568 1414
rect 5092 800 5120 3334
rect 5184 3126 5212 4134
rect 5276 3534 5304 4966
rect 5368 3738 5396 6886
rect 6104 5710 6132 7142
rect 6288 6662 6316 11104
rect 6368 11144 6420 11150
rect 6472 11132 6500 11494
rect 6420 11104 6500 11132
rect 6368 11086 6420 11092
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9654 6408 9930
rect 6472 9926 6500 11104
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 7410 6408 8366
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6380 7206 6408 7346
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6472 6914 6500 9862
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7410 6684 7686
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6380 6886 6500 6914
rect 6748 6914 6776 11766
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11280 6880 11286
rect 6828 11222 6880 11228
rect 6840 10962 6868 11222
rect 6932 11150 6960 11630
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6840 10934 6960 10962
rect 6932 10606 6960 10934
rect 7024 10810 7052 11154
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7116 10674 7144 11834
rect 7208 11762 7236 12056
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11286 7236 11698
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7208 10062 7236 11086
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8566 7052 8774
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7478 6960 7686
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7208 6914 7236 9998
rect 6748 6886 6868 6914
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 4622 6132 5646
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5448 4208 5500 4214
rect 5552 4185 5580 4558
rect 5448 4150 5500 4156
rect 5538 4176 5594 4185
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5460 2990 5488 4150
rect 5538 4111 5540 4120
rect 5592 4111 5594 4120
rect 5540 4082 5592 4088
rect 5552 3534 5580 4082
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 2854 5488 2926
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5552 800 5580 2518
rect 6288 2514 6316 6598
rect 6276 2508 6328 2514
rect 6276 2450 6328 2456
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6012 800 6040 2246
rect 6380 2106 6408 6886
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4282 6684 4490
rect 6748 4282 6776 4966
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6458 3496 6514 3505
rect 6458 3431 6514 3440
rect 6472 3398 6500 3431
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6564 3058 6592 4082
rect 6748 4078 6776 4218
rect 6840 4146 6868 6886
rect 7116 6886 7236 6914
rect 7116 6798 7144 6886
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5370 7144 6598
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6932 4622 6960 5170
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7116 4486 7144 5170
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6656 3738 6684 4014
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3670 6776 3878
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6748 2938 6776 3470
rect 6840 3126 6868 4082
rect 6918 3768 6974 3777
rect 7208 3738 7236 5510
rect 7300 5370 7328 19110
rect 7392 18970 7420 21966
rect 7472 21888 7524 21894
rect 7472 21830 7524 21836
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7392 18766 7420 18906
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7484 18612 7512 21830
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 7576 20874 7604 21626
rect 7668 21078 7696 23190
rect 7840 23044 7892 23050
rect 7840 22986 7892 22992
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7760 21894 7788 22510
rect 7852 22094 7880 22986
rect 7852 22066 8156 22094
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7760 21690 7788 21830
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 8128 21554 8156 22066
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21554 8248 21898
rect 7748 21548 7800 21554
rect 8116 21548 8168 21554
rect 7800 21508 7880 21536
rect 7748 21490 7800 21496
rect 7852 21350 7880 21508
rect 8116 21490 8168 21496
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7748 21344 7800 21350
rect 7748 21286 7800 21292
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7760 21146 7788 21286
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7840 21140 7892 21146
rect 7840 21082 7892 21088
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7392 18584 7512 18612
rect 7392 13530 7420 18584
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 16998 7512 17478
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7576 15026 7604 20810
rect 7668 20262 7696 21014
rect 7852 20942 7880 21082
rect 8036 21026 8064 21422
rect 7944 20998 8064 21026
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7760 20398 7788 20878
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7852 19514 7880 20402
rect 7944 19854 7972 20998
rect 8024 20912 8076 20918
rect 8024 20854 8076 20860
rect 8036 20602 8064 20854
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 8128 20534 8156 21490
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7576 13394 7604 14758
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7668 13326 7696 14418
rect 7760 14414 7788 18838
rect 7944 18766 7972 19654
rect 8036 19174 8064 19722
rect 8128 19242 8156 19722
rect 8220 19446 8248 21286
rect 9324 21078 9352 26318
rect 9600 25294 9628 27406
rect 10508 27396 10560 27402
rect 10508 27338 10560 27344
rect 10520 27130 10548 27338
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 10888 27130 10916 27270
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10980 26382 11008 26930
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9588 23520 9640 23526
rect 9640 23468 9720 23474
rect 9588 23462 9720 23468
rect 9600 23446 9720 23462
rect 9692 22098 9720 23446
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8312 19378 8340 19994
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 8128 18612 8156 19178
rect 8680 18766 8708 20742
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8864 18834 8892 20402
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 7944 18584 8156 18612
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 17202 7880 18226
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 15910 7880 17138
rect 7944 15910 7972 18584
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7760 14006 7788 14350
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7576 12850 7604 13194
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7380 12164 7432 12170
rect 7380 12106 7432 12112
rect 7392 11150 7420 12106
rect 7484 11830 7512 12310
rect 7668 11830 7696 13262
rect 7760 12986 7788 13942
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 12238 7788 12718
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11218 7604 11698
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10674 7420 11086
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7760 10606 7788 12174
rect 7852 11694 7880 13874
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 9382 7512 9522
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 8974 7512 9318
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8634 7420 8774
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7484 8498 7512 8910
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 7886 7512 8434
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7484 4826 7512 6734
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 6918 3703 6974 3712
rect 7196 3732 7248 3738
rect 6932 3670 6960 3703
rect 7196 3674 7248 3680
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6748 2922 7328 2938
rect 6748 2916 7340 2922
rect 6748 2910 7288 2916
rect 7288 2858 7340 2864
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6368 2100 6420 2106
rect 6368 2042 6420 2048
rect 6472 870 6592 898
rect 6472 800 6500 870
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6564 762 6592 870
rect 6748 762 6776 2246
rect 7116 1494 7144 2382
rect 7104 1488 7156 1494
rect 7104 1430 7156 1436
rect 7484 800 7512 3470
rect 7576 3058 7604 10406
rect 7760 5794 7788 10406
rect 7852 10130 7880 10610
rect 7944 10538 7972 13398
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7852 6730 7880 10066
rect 8036 6934 8064 18022
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8128 16046 8156 16458
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 5914 7880 6666
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7760 5766 8064 5794
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7944 4826 7972 5578
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7760 3738 7788 4558
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3534 7880 4422
rect 7944 4282 7972 4558
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8036 4078 8064 5766
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8128 3942 8156 15846
rect 8220 15162 8248 18634
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 14346 8248 15098
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8220 13938 8248 14282
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8588 13462 8616 14826
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8588 12850 8616 13398
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8680 11558 8708 18702
rect 8864 15026 8892 18770
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17882 8984 18226
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 9310 17776 9366 17785
rect 9310 17711 9366 17720
rect 9128 17672 9180 17678
rect 9126 17640 9128 17649
rect 9220 17672 9272 17678
rect 9180 17640 9182 17649
rect 9220 17614 9272 17620
rect 9126 17575 9182 17584
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17202 9168 17478
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8956 16794 8984 17138
rect 9126 17096 9182 17105
rect 9126 17031 9182 17040
rect 9140 16998 9168 17031
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 9140 16454 9168 16934
rect 9232 16658 9260 17614
rect 9324 17610 9352 17711
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 8852 15020 8904 15026
rect 8772 14980 8852 15008
rect 8772 11898 8800 14980
rect 8852 14962 8904 14968
rect 9416 13274 9444 19314
rect 9494 17776 9550 17785
rect 9494 17711 9496 17720
rect 9548 17711 9550 17720
rect 9496 17682 9548 17688
rect 9494 17640 9550 17649
rect 9494 17575 9550 17584
rect 9508 17542 9536 17575
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9508 14346 9536 15098
rect 9600 14618 9628 20198
rect 9692 18426 9720 20266
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9692 17678 9720 18362
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9784 14521 9812 24754
rect 9876 20330 9904 25094
rect 10060 24886 10088 25094
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 10152 24818 10180 26318
rect 12084 26234 12112 36722
rect 12900 30796 12952 30802
rect 12900 30738 12952 30744
rect 12912 29306 12940 30738
rect 12900 29300 12952 29306
rect 12900 29242 12952 29248
rect 12348 29232 12400 29238
rect 12348 29174 12400 29180
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 12176 28762 12204 29106
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 12360 27538 12388 29174
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12360 26994 12388 27474
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12360 26466 12388 26930
rect 12636 26586 12664 28494
rect 12912 28490 12940 29242
rect 12900 28484 12952 28490
rect 12900 28426 12952 28432
rect 13176 27056 13228 27062
rect 13176 26998 13228 27004
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12360 26438 12480 26466
rect 12348 26308 12400 26314
rect 12348 26250 12400 26256
rect 12084 26206 12204 26234
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10244 24954 10272 25162
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10152 24274 10180 24754
rect 10600 24744 10652 24750
rect 10600 24686 10652 24692
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10336 24342 10364 24618
rect 10324 24336 10376 24342
rect 10324 24278 10376 24284
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10152 23798 10180 24210
rect 10336 24206 10364 24278
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 10152 23610 10180 23734
rect 10060 23582 10180 23610
rect 10244 23594 10272 24142
rect 10232 23588 10284 23594
rect 10060 23186 10088 23582
rect 10232 23530 10284 23536
rect 10244 23474 10272 23530
rect 10152 23446 10272 23474
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10152 23118 10180 23446
rect 10336 23254 10364 24142
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 10428 23322 10456 23666
rect 10520 23497 10548 24142
rect 10612 24138 10640 24686
rect 11072 24410 11100 25162
rect 12176 25158 12204 26206
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 12176 24138 12204 25094
rect 10600 24132 10652 24138
rect 10600 24074 10652 24080
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 10506 23488 10562 23497
rect 10506 23423 10562 23432
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9968 14822 9996 23054
rect 10612 23050 10640 24074
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 12084 23118 12112 23666
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10600 23044 10652 23050
rect 10600 22986 10652 22992
rect 10336 22438 10364 22986
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 10244 19922 10272 22034
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 18714 10272 19858
rect 10152 18686 10272 18714
rect 10152 18358 10180 18686
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 14890 10180 17138
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9770 14512 9826 14521
rect 9770 14447 9826 14456
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9508 13394 9536 14282
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9600 13326 9628 14214
rect 9588 13320 9640 13326
rect 9416 13246 9536 13274
rect 9588 13262 9640 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12306 9444 13126
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9036 12232 9088 12238
rect 9220 12232 9272 12238
rect 9088 12192 9220 12220
rect 9036 12174 9088 12180
rect 9220 12174 9272 12180
rect 9416 12102 9444 12242
rect 9508 12238 9536 13246
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9968 12889 9996 12922
rect 9954 12880 10010 12889
rect 9954 12815 10010 12824
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 9680 12640 9732 12646
rect 9678 12608 9680 12617
rect 9732 12608 9734 12617
rect 9678 12543 9734 12552
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 6186 8340 8366
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8036 3534 8064 3878
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8312 3194 8340 5306
rect 8404 4146 8432 9318
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8404 3058 8432 3130
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 7944 800 7972 2246
rect 8496 800 8524 2246
rect 8588 1086 8616 4082
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 3058 8708 3334
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8772 2378 8800 11698
rect 8864 9586 8892 12038
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 9692 9466 9720 12038
rect 10152 11762 10180 12718
rect 10244 12374 10272 18566
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10230 12200 10286 12209
rect 10230 12135 10286 12144
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9508 9438 9720 9466
rect 9508 9178 9536 9438
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9508 8498 9536 8978
rect 9692 8974 9720 9318
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9600 7206 9628 8910
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 6254 9628 7142
rect 9692 7002 9720 7346
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6882 9812 11222
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9968 9586 9996 11018
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9876 8634 9904 9522
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9968 8514 9996 9318
rect 9876 8486 9996 8514
rect 9876 7886 9904 8486
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9692 6866 9812 6882
rect 9680 6860 9812 6866
rect 9732 6854 9812 6860
rect 9680 6802 9732 6808
rect 9876 6474 9904 7822
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9968 6934 9996 7754
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9968 6662 9996 6870
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9876 6446 9996 6474
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 2514 8892 6054
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 3505 9168 3674
rect 9324 3670 9352 4150
rect 9312 3664 9364 3670
rect 9218 3632 9274 3641
rect 9312 3606 9364 3612
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9218 3567 9220 3576
rect 9272 3567 9274 3576
rect 9220 3538 9272 3544
rect 9126 3496 9182 3505
rect 9126 3431 9182 3440
rect 9416 3126 9444 3606
rect 9508 3534 9536 5578
rect 9600 5098 9628 6190
rect 9876 5914 9904 6258
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9600 4146 9628 4694
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9600 3194 9628 4082
rect 9784 3942 9812 4558
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9692 3534 9720 3878
rect 9784 3534 9812 3878
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9968 3058 9996 6446
rect 10060 5302 10088 11018
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10152 5710 10180 10134
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10060 4826 10088 5238
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10152 4690 10180 5034
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10152 2990 10180 3946
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8576 1080 8628 1086
rect 8576 1022 8628 1028
rect 8956 870 9076 898
rect 8956 800 8984 870
rect 6564 734 6776 762
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9048 762 9076 870
rect 9232 762 9260 2246
rect 9416 800 9444 2518
rect 9784 2446 9812 2790
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10244 1698 10272 12135
rect 10336 5710 10364 22374
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20602 10548 20878
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 12102 10456 20334
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10520 15706 10548 16050
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10612 15570 10640 20266
rect 10704 19854 10732 20742
rect 11072 20602 11100 20742
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 20058 11836 20402
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 11808 19446 11836 19994
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 13938 10548 14350
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13462 10548 13874
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12850 10548 13126
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10506 12744 10562 12753
rect 10506 12679 10562 12688
rect 10520 12238 10548 12679
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10416 12096 10468 12102
rect 10612 12084 10640 15506
rect 10704 12850 10732 18634
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 10874 16688 10930 16697
rect 10874 16623 10876 16632
rect 10928 16623 10930 16632
rect 10876 16594 10928 16600
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 16250 10824 16458
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16250 10916 16390
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15502 10916 15846
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10796 14414 10824 14554
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 14278 10824 14350
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10612 12056 10732 12084
rect 10416 12038 10468 12044
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 6914 10456 11494
rect 10520 10742 10548 11698
rect 10612 11354 10640 11698
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10520 9382 10548 10474
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10612 9450 10640 9590
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8634 10548 8774
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10612 7886 10640 9386
rect 10704 8430 10732 12056
rect 10796 11150 10824 12310
rect 10888 12238 10916 12786
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10796 6914 10824 10950
rect 10888 10538 10916 12174
rect 10980 10826 11008 12582
rect 11072 11286 11100 15302
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11164 11014 11192 14758
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10980 10810 11100 10826
rect 10980 10804 11112 10810
rect 10980 10798 11060 10804
rect 11060 10746 11112 10752
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10428 6886 10548 6914
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10336 5302 10364 5646
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10520 5234 10548 6886
rect 10704 6886 10824 6914
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4622 10456 4966
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10232 1692 10284 1698
rect 10232 1634 10284 1640
rect 10428 800 10456 4082
rect 10612 4010 10640 6258
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10600 3528 10652 3534
rect 10598 3496 10600 3505
rect 10652 3496 10654 3505
rect 10598 3431 10654 3440
rect 10704 1630 10732 6886
rect 10888 6390 10916 9862
rect 10980 9654 11008 10678
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 9178 11008 9590
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11440 7886 11468 18158
rect 11900 16046 11928 22918
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 11992 16726 12020 17002
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11624 14006 11652 14486
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 6798 11100 7686
rect 11440 7274 11468 7822
rect 11532 7750 11560 13942
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11624 11286 11652 12242
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11624 10674 11652 11222
rect 11716 10674 11744 13670
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11808 11354 11836 11698
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10062 11652 10406
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11716 10062 11744 10202
rect 11900 10062 11928 15982
rect 12084 15162 12112 23054
rect 12360 22982 12388 26250
rect 12452 25906 12480 26438
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12452 25294 12480 25842
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12452 24290 12480 25230
rect 12452 24274 12572 24290
rect 12452 24268 12584 24274
rect 12452 24262 12532 24268
rect 12452 23662 12480 24262
rect 12532 24210 12584 24216
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20534 12480 20810
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12360 18290 12388 19314
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12544 18766 12572 18838
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12728 18630 12756 24142
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17202 12204 17478
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12268 17066 12296 17614
rect 12360 17202 12388 18226
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12268 16794 12296 17002
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13938 12020 14214
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 10266 12020 11698
rect 12084 11150 12112 15098
rect 12176 14958 12204 15098
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12360 13734 12388 17138
rect 12636 16454 12664 17750
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 16998 12756 17614
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14074 12480 14894
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12636 13530 12664 14962
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12617 12572 12854
rect 12530 12608 12586 12617
rect 12530 12543 12586 12552
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11900 9722 11928 9998
rect 12360 9722 12388 11086
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11716 9178 11744 9454
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 12360 8974 12388 9658
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11716 8634 11744 8842
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11532 6914 11560 7686
rect 12544 7206 12572 11698
rect 12636 11694 12664 13466
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 7546 12756 8434
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 11348 6886 11560 6914
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 11072 5778 11100 6734
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10796 3398 10824 3946
rect 11348 3942 11376 6886
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10888 3641 10916 3674
rect 10874 3632 10930 3641
rect 10874 3567 10930 3576
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10692 1624 10744 1630
rect 10692 1566 10744 1572
rect 10888 800 10916 3402
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10980 3058 11008 3334
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11900 2650 11928 6190
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12452 3777 12480 5782
rect 12544 4214 12572 7142
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12438 3768 12494 3777
rect 12438 3703 12494 3712
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 12268 2446 12296 2790
rect 12820 2774 12848 24074
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12912 22030 12940 22986
rect 13004 22098 13032 23462
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12912 20058 12940 20470
rect 13096 20262 13124 22646
rect 13188 22094 13216 26998
rect 13280 24206 13308 38898
rect 14464 38344 14516 38350
rect 14464 38286 14516 38292
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13648 24206 13676 24754
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13280 23746 13308 24142
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13372 23866 13400 24006
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13556 23798 13584 24006
rect 13544 23792 13596 23798
rect 13280 23718 13492 23746
rect 13544 23734 13596 23740
rect 13464 23526 13492 23718
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13648 23254 13676 24142
rect 13636 23248 13688 23254
rect 13636 23190 13688 23196
rect 13740 22438 13768 28358
rect 14476 27130 14504 38286
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 15476 31952 15528 31958
rect 15476 31894 15528 31900
rect 15488 29306 15516 31894
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14752 28762 14780 29106
rect 14740 28756 14792 28762
rect 14740 28698 14792 28704
rect 15488 28490 15516 29242
rect 15476 28484 15528 28490
rect 15476 28426 15528 28432
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14004 26444 14056 26450
rect 14004 26386 14056 26392
rect 14016 24614 14044 26386
rect 14476 26382 14504 27066
rect 15304 26994 15332 27474
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 14752 26586 14780 26930
rect 14740 26580 14792 26586
rect 14740 26522 14792 26528
rect 15304 26450 15332 26930
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14096 26240 14148 26246
rect 14096 26182 14148 26188
rect 14108 25294 14136 26182
rect 14384 25974 14412 26250
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14384 25226 14412 25910
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25294 14504 25638
rect 14568 25294 14596 26318
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 16212 26308 16264 26314
rect 16212 26250 16264 26256
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14752 25430 14780 25842
rect 14740 25424 14792 25430
rect 14740 25366 14792 25372
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14384 24138 14412 25162
rect 14568 24818 14596 25230
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14384 23798 14412 24074
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14844 23322 14872 23734
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14844 22642 14872 23054
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13188 22066 13584 22094
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13188 20074 13216 20470
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13096 20046 13216 20074
rect 12912 19378 12940 19994
rect 13096 19854 13124 20046
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 5642 12940 18566
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 16726 13032 17546
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13096 16522 13124 19790
rect 13372 19378 13400 20946
rect 13556 19514 13584 22066
rect 14188 22024 14240 22030
rect 14292 22012 14320 22510
rect 14240 21984 14320 22012
rect 14188 21966 14240 21972
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13832 21690 13860 21898
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 14292 21554 14320 21984
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14568 21146 14596 21490
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13740 19922 13768 20810
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13648 19378 13676 19790
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17202 13400 17614
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 16726 13400 17138
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13096 13870 13124 16458
rect 13372 15026 13400 16662
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13280 14618 13308 14758
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13096 12850 13124 13806
rect 13280 13394 13308 13806
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13280 12782 13308 13330
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13372 9586 13400 14962
rect 13464 13870 13492 19178
rect 14016 19145 14044 19246
rect 14002 19136 14058 19145
rect 14002 19071 14058 19080
rect 14464 18148 14516 18154
rect 14464 18090 14516 18096
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 16697 13860 17614
rect 14476 16998 14504 18090
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 13818 16688 13874 16697
rect 13818 16623 13874 16632
rect 13832 16046 13860 16623
rect 13924 16289 13952 16934
rect 13910 16280 13966 16289
rect 13910 16215 13966 16224
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13556 14074 13584 15030
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13464 12714 13492 13806
rect 13832 13734 13860 14758
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13924 13190 13952 16215
rect 14476 16114 14504 16934
rect 14568 16522 14596 21082
rect 14844 20330 14872 22578
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14646 16824 14702 16833
rect 14752 16794 14780 17478
rect 14936 17218 14964 26250
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15212 25906 15240 26182
rect 16224 26042 16252 26250
rect 16212 26036 16264 26042
rect 16212 25978 16264 25984
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 15016 25152 15068 25158
rect 15016 25094 15068 25100
rect 14844 17190 14964 17218
rect 14646 16759 14648 16768
rect 14700 16759 14702 16768
rect 14740 16788 14792 16794
rect 14648 16730 14700 16736
rect 14740 16730 14792 16736
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 14482 14412 15982
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13452 12708 13504 12714
rect 13452 12650 13504 12656
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11830 13584 12038
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13004 8362 13032 9454
rect 13372 8498 13400 9522
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 13096 7954 13124 8298
rect 13464 8294 13492 8502
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13188 7546 13216 7822
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13280 7002 13308 7822
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 5846 13124 6734
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 6322 13308 6666
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 13556 4554 13584 9318
rect 13648 4622 13676 12582
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 11082 13768 11766
rect 13832 11694 13860 11834
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13924 9518 13952 13126
rect 14384 12714 14412 14418
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14384 12434 14412 12650
rect 14292 12406 14412 12434
rect 14292 12238 14320 12406
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13740 7002 13768 7958
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13740 6798 13768 6938
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13832 5710 13860 8434
rect 13924 7410 13952 8978
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3602 13032 4082
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13004 3058 13032 3538
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12728 2746 12848 2774
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 11336 2304 11388 2310
rect 11336 2246 11388 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11348 800 11376 2246
rect 11900 800 11928 2246
rect 12360 800 12388 2518
rect 12728 1766 12756 2746
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13004 2038 13032 2382
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12716 1760 12768 1766
rect 12716 1702 12768 1708
rect 13372 800 13400 3402
rect 13832 800 13860 4150
rect 13924 3602 13952 7346
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 3058 13952 3538
rect 14016 3534 14044 10542
rect 14108 7886 14136 10678
rect 14292 10674 14320 12174
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14384 10742 14412 11018
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14660 10266 14688 16730
rect 14844 12434 14872 17190
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15706 14964 16050
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 15028 15586 15056 25094
rect 15212 23730 15240 25842
rect 15948 24818 15976 25842
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15488 24274 15516 24686
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15212 23526 15240 23666
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15488 23186 15516 24210
rect 15672 23730 15700 24754
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15856 23866 15884 24074
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 15120 19718 15148 20266
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15212 18222 15240 21830
rect 15488 21622 15516 21830
rect 15476 21616 15528 21622
rect 15476 21558 15528 21564
rect 15568 21616 15620 21622
rect 15568 21558 15620 21564
rect 15580 20806 15608 21558
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15672 21146 15700 21422
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15672 20618 15700 20946
rect 15580 20590 15700 20618
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15384 19848 15436 19854
rect 15488 19802 15516 20334
rect 15580 20330 15608 20590
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15580 19922 15608 20266
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 15436 19796 15516 19802
rect 15384 19790 15516 19796
rect 15396 19774 15516 19790
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15304 19378 15332 19654
rect 15396 19514 15424 19654
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15488 18290 15516 19774
rect 15568 19780 15620 19786
rect 15620 19740 15700 19768
rect 15568 19722 15620 19728
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15580 18426 15608 18634
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 17338 15148 17478
rect 15304 17338 15332 17546
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15396 16998 15424 17138
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15396 16182 15424 16458
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 14752 12406 14872 12434
rect 14936 15558 15056 15586
rect 15290 15600 15346 15609
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14292 9586 14320 10202
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14752 9602 14780 12406
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14844 9722 14872 9930
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8974 14412 9318
rect 14568 8974 14596 9590
rect 14752 9574 14872 9602
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14660 9042 14688 9454
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14372 8968 14424 8974
rect 14292 8928 14372 8956
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8498 14228 8774
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6798 14136 7210
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14200 6662 14228 7822
rect 14292 7478 14320 8928
rect 14372 8910 14424 8916
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14568 8786 14596 8910
rect 14568 8758 14688 8786
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14568 8430 14596 8502
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7954 14596 8366
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14292 6118 14320 6734
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14476 5710 14504 7346
rect 14660 7342 14688 8758
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14660 6798 14688 6938
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14752 6662 14780 8434
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5302 14136 5510
rect 14476 5370 14504 5646
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14844 2922 14872 9574
rect 14936 7970 14964 15558
rect 15290 15535 15292 15544
rect 15344 15535 15346 15544
rect 15292 15506 15344 15512
rect 15108 15496 15160 15502
rect 15160 15456 15240 15484
rect 15108 15438 15160 15444
rect 15212 14958 15240 15456
rect 15200 14952 15252 14958
rect 15304 14940 15332 15506
rect 15396 15434 15424 16118
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15384 14952 15436 14958
rect 15304 14912 15384 14940
rect 15200 14894 15252 14900
rect 15384 14894 15436 14900
rect 15212 14822 15240 14894
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15028 14414 15056 14758
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 11898 15148 12106
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15212 11744 15240 14758
rect 15396 14498 15424 14894
rect 15488 14618 15516 18226
rect 15672 17882 15700 19740
rect 15764 18630 15792 23462
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 15856 20942 15884 21354
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 15856 19718 15884 20878
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15948 19854 15976 19994
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15856 18902 15884 19178
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15948 18630 15976 19450
rect 15752 18624 15804 18630
rect 15936 18624 15988 18630
rect 15804 18572 15884 18578
rect 15752 18566 15884 18572
rect 15936 18566 15988 18572
rect 15764 18550 15884 18566
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15672 17338 15700 17818
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15764 15978 15792 18294
rect 15752 15972 15804 15978
rect 15752 15914 15804 15920
rect 15764 15434 15792 15914
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15396 14470 15792 14498
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 14074 15700 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15304 12102 15332 12854
rect 15488 12646 15516 14010
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11756 15344 11762
rect 15212 11716 15292 11744
rect 15212 11218 15240 11716
rect 15292 11698 15344 11704
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15292 11144 15344 11150
rect 15396 11132 15424 11834
rect 15488 11354 15516 12582
rect 15672 11762 15700 12582
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15764 11694 15792 14470
rect 15856 13870 15884 18550
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15948 12170 15976 18566
rect 16040 14618 16068 20878
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 16132 19446 16160 19722
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16132 18290 16160 19246
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16224 17882 16252 21286
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16132 17338 16160 17614
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16132 14618 16160 15642
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16040 14346 16068 14554
rect 16316 14498 16344 15302
rect 16132 14470 16344 14498
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16132 13190 16160 14470
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12918 16160 13126
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15764 11150 15792 11630
rect 15344 11104 15424 11132
rect 15292 11086 15344 11092
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10742 15056 10950
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15212 9994 15240 10678
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14936 7942 15056 7970
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14936 3670 14964 6802
rect 15028 4214 15056 7942
rect 15212 7410 15240 9930
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 15120 3194 15148 4082
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15120 2446 15148 2790
rect 15212 2553 15240 2790
rect 15198 2544 15254 2553
rect 15304 2514 15332 6394
rect 15396 5234 15424 11104
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8560 15712 8566
rect 15488 8508 15660 8514
rect 15488 8502 15712 8508
rect 15488 8486 15700 8502
rect 15764 8498 15792 8774
rect 15752 8492 15804 8498
rect 15488 8430 15516 8486
rect 15752 8434 15804 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15948 7954 15976 12106
rect 16132 11082 16160 12854
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16040 10470 16068 11018
rect 16224 10962 16252 13806
rect 16316 12714 16344 13942
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 16408 12434 16436 25774
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16132 10934 16252 10962
rect 16316 12406 16436 12434
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 16132 7818 16160 10934
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 7818 16252 8434
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16132 7002 16160 7210
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16132 6798 16160 6938
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16224 6322 16252 6870
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 3602 15516 4966
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15488 3398 15516 3538
rect 15764 3534 15792 4422
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15396 3058 15424 3334
rect 16040 3058 16068 3878
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15198 2479 15254 2488
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 14292 800 14320 2246
rect 14844 800 14872 2246
rect 15396 1170 15424 2246
rect 15304 1142 15424 1170
rect 15304 800 15332 1142
rect 16224 800 16252 4082
rect 16316 1970 16344 12406
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 10742 16436 12038
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16396 10532 16448 10538
rect 16396 10474 16448 10480
rect 16408 5710 16436 10474
rect 16396 5704 16448 5710
rect 16396 5646 16448 5652
rect 16408 4690 16436 5646
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16500 2774 16528 23598
rect 16592 21690 16620 28358
rect 17052 28218 17080 32846
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17040 28212 17092 28218
rect 17040 28154 17092 28160
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16684 27470 16712 27814
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 16776 25974 16804 26522
rect 16764 25968 16816 25974
rect 16764 25910 16816 25916
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16776 22778 16804 22986
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16592 20466 16620 21490
rect 16868 21146 16896 28018
rect 17052 27674 17080 28154
rect 17144 28082 17172 28494
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 17328 26994 17356 28494
rect 18052 28484 18104 28490
rect 18052 28426 18104 28432
rect 18064 28218 18092 28426
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 18708 28150 18736 28358
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 18696 28144 18748 28150
rect 18696 28086 18748 28092
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18156 26586 18184 26930
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23798 16988 24006
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22710 17448 22918
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 16948 22636 17000 22642
rect 17000 22596 17080 22624
rect 16948 22578 17000 22584
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16960 20534 16988 21422
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 17052 19514 17080 22596
rect 18248 22098 18276 28018
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18604 26784 18656 26790
rect 18604 26726 18656 26732
rect 18616 26382 18644 26726
rect 18708 26382 18736 27950
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 24410 18368 24754
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17420 21010 17448 21286
rect 17604 21146 17632 21490
rect 17880 21486 17908 21830
rect 18432 21690 18460 26318
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 24138 18644 24550
rect 18892 24274 18920 24686
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18708 23526 18736 24142
rect 19064 24132 19116 24138
rect 19064 24074 19116 24080
rect 19076 23866 19104 24074
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18708 22778 18736 23462
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 19156 22636 19208 22642
rect 19524 22636 19576 22642
rect 19156 22578 19208 22584
rect 19444 22596 19524 22624
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18616 22166 18644 22510
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18616 21622 18644 22102
rect 18708 22030 18736 22510
rect 18880 22160 18932 22166
rect 18880 22102 18932 22108
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17604 21010 17632 21082
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17696 20942 17724 21422
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17144 19378 17172 20402
rect 17512 20058 17540 20878
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17696 19854 17724 20878
rect 17880 20806 17908 21422
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17880 20398 17908 20742
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17972 20330 18000 21490
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18156 20874 18184 21422
rect 18616 21146 18644 21558
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18708 20942 18736 21966
rect 18800 21554 18828 21966
rect 18892 21554 18920 22102
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18984 21350 19012 22578
rect 19168 21486 19196 22578
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22234 19288 22374
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19444 22137 19472 22596
rect 19524 22578 19576 22584
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19430 22128 19486 22137
rect 19536 22098 19564 22442
rect 19812 22438 19840 22578
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19812 22098 19840 22374
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19430 22063 19486 22072
rect 19524 22092 19576 22098
rect 19444 22030 19472 22063
rect 19524 22034 19576 22040
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 19352 21146 19380 21422
rect 19444 21185 19472 21966
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19430 21176 19486 21185
rect 19340 21140 19392 21146
rect 19430 21111 19486 21120
rect 19340 21082 19392 21088
rect 19616 21072 19668 21078
rect 19668 21032 19748 21060
rect 19616 21014 19668 21020
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 19294 20936 19346 20942
rect 19294 20878 19346 20884
rect 19430 20904 19486 20913
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 18052 20460 18104 20466
rect 18156 20448 18184 20810
rect 18104 20420 18184 20448
rect 18052 20402 18104 20408
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18432 19922 18460 20334
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17420 19446 17448 19790
rect 17408 19440 17460 19446
rect 17408 19382 17460 19388
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17144 18970 17172 19314
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16592 14618 16620 14962
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16684 12238 16712 18226
rect 17052 17116 17080 18838
rect 17316 18760 17368 18766
rect 17420 18748 17448 19382
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 17368 18720 17448 18748
rect 17316 18702 17368 18708
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17236 18290 17264 18362
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17972 18222 18000 18838
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17144 17610 17172 18158
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17132 17128 17184 17134
rect 17052 17088 17132 17116
rect 17132 17070 17184 17076
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17052 16046 17080 16730
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16592 10130 16620 10610
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16684 9586 16712 12174
rect 17144 10674 17172 17070
rect 17512 16153 17540 17070
rect 17498 16144 17554 16153
rect 17498 16079 17500 16088
rect 17552 16079 17554 16088
rect 17500 16050 17552 16056
rect 17316 16040 17368 16046
rect 18064 15994 18092 19110
rect 18340 18426 18368 19314
rect 18432 19174 18460 19858
rect 19168 19310 19196 20810
rect 19306 20602 19334 20878
rect 19536 20890 19564 20946
rect 19720 20942 19748 21032
rect 19708 20936 19760 20942
rect 19614 20904 19670 20913
rect 19536 20862 19614 20890
rect 19430 20839 19486 20848
rect 19708 20878 19760 20884
rect 19614 20839 19670 20848
rect 19294 20596 19346 20602
rect 19444 20584 19472 20839
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19444 20556 19840 20584
rect 19294 20538 19346 20544
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19260 19378 19288 20402
rect 19352 20369 19380 20402
rect 19524 20392 19576 20398
rect 19338 20360 19394 20369
rect 19524 20334 19576 20340
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19338 20295 19394 20304
rect 19536 20233 19564 20334
rect 19522 20224 19578 20233
rect 19522 20159 19578 20168
rect 19720 19922 19748 20334
rect 19812 19922 19840 20556
rect 19892 20392 19944 20398
rect 19890 20360 19892 20369
rect 19944 20360 19946 20369
rect 19890 20295 19946 20304
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19892 19848 19944 19854
rect 19996 19836 20024 22102
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20088 20398 20116 21422
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19944 19808 20024 19836
rect 19892 19790 19944 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 19154 19136 19210 19145
rect 19154 19071 19210 19080
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18328 18420 18380 18426
rect 18380 18380 18552 18408
rect 18328 18362 18380 18368
rect 18340 18297 18368 18362
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 18086 18184 18158
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18144 17536 18196 17542
rect 18248 17524 18276 17818
rect 18340 17678 18368 18022
rect 18524 17746 18552 18380
rect 18616 18290 18644 18770
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 19076 18154 19104 18226
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18616 17746 18828 17762
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18616 17740 18840 17746
rect 18616 17734 18788 17740
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18196 17496 18276 17524
rect 18144 17478 18196 17484
rect 18432 17270 18460 17614
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16969 18552 17138
rect 18616 17134 18644 17734
rect 18788 17682 18840 17688
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18510 16960 18566 16969
rect 18510 16895 18566 16904
rect 18616 16833 18644 17070
rect 18602 16824 18658 16833
rect 18602 16759 18658 16768
rect 18708 16590 18736 17614
rect 19076 17202 19104 18090
rect 19168 17202 19196 19071
rect 19536 18970 19564 19246
rect 19720 19009 19748 19246
rect 19904 19174 19932 19246
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19706 19000 19762 19009
rect 19524 18964 19576 18970
rect 19904 18970 19932 19110
rect 19706 18935 19762 18944
rect 19892 18964 19944 18970
rect 19524 18906 19576 18912
rect 19892 18906 19944 18912
rect 19708 18760 19760 18766
rect 19996 18748 20024 19808
rect 20088 19174 20116 20334
rect 20180 19786 20208 20538
rect 20272 20233 20300 24006
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20364 22234 20392 22714
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20444 22024 20496 22030
rect 20350 21992 20406 22001
rect 20444 21966 20496 21972
rect 20350 21927 20352 21936
rect 20404 21927 20406 21936
rect 20352 21898 20404 21904
rect 20456 21690 20484 21966
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20352 20256 20404 20262
rect 20258 20224 20314 20233
rect 20352 20198 20404 20204
rect 20258 20159 20314 20168
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20272 18834 20300 19858
rect 20364 19786 20392 20198
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20548 18970 20576 23802
rect 20640 23798 20668 24006
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22574 21680 23054
rect 21732 22976 21784 22982
rect 21732 22918 21784 22924
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20626 22128 20682 22137
rect 20626 22063 20628 22072
rect 20680 22063 20682 22072
rect 20628 22034 20680 22040
rect 20824 22030 20852 22170
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 21652 20942 21680 22510
rect 21744 22506 21772 22918
rect 21732 22500 21784 22506
rect 21732 22442 21784 22448
rect 21744 21962 21772 22442
rect 21928 22094 21956 32166
rect 25504 27396 25556 27402
rect 25504 27338 25556 27344
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 21836 22066 21956 22094
rect 21732 21956 21784 21962
rect 21732 21898 21784 21904
rect 21640 20936 21692 20942
rect 20626 20904 20682 20913
rect 21640 20878 21692 20884
rect 20626 20839 20682 20848
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 19760 18720 20024 18748
rect 19708 18702 19760 18708
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19260 18222 19288 18634
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19996 18290 20024 18720
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19996 17678 20024 18226
rect 20272 18204 20300 18770
rect 20640 18222 20668 20839
rect 21652 19854 21680 20878
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 21744 20262 21772 20470
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21652 19378 21680 19790
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 18426 20760 18702
rect 20824 18426 20852 19178
rect 20916 18766 20944 19246
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18766 21036 19110
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20444 18216 20496 18222
rect 20272 18176 20444 18204
rect 20444 18158 20496 18164
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21560 17814 21588 18022
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 20628 17536 20680 17542
rect 20626 17504 20628 17513
rect 20680 17504 20682 17513
rect 19574 17436 19882 17456
rect 20626 17439 20682 17448
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 18878 16960 18934 16969
rect 18878 16895 18934 16904
rect 18892 16726 18920 16895
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18340 16250 18368 16526
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18432 16114 18460 16458
rect 18708 16153 18736 16526
rect 18786 16280 18842 16289
rect 18786 16215 18842 16224
rect 18800 16182 18828 16215
rect 18788 16176 18840 16182
rect 18694 16144 18750 16153
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18420 16108 18472 16114
rect 18788 16118 18840 16124
rect 19076 16114 19104 17138
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 21652 16182 21680 17614
rect 21730 17096 21786 17105
rect 21730 17031 21786 17040
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 18694 16079 18696 16088
rect 18420 16050 18472 16056
rect 18748 16079 18750 16088
rect 19064 16108 19116 16114
rect 18696 16050 18748 16056
rect 19064 16050 19116 16056
rect 17316 15982 17368 15988
rect 17328 13802 17356 15982
rect 17972 15966 18092 15994
rect 17972 15858 18000 15966
rect 17880 15830 18000 15858
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17880 15042 17908 15830
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 15162 18000 15642
rect 18064 15570 18092 15846
rect 18248 15706 18276 16050
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18064 15178 18092 15506
rect 18340 15502 18368 15642
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 17960 15156 18012 15162
rect 18064 15150 18276 15178
rect 17960 15098 18012 15104
rect 17880 15014 18000 15042
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17236 13530 17264 13738
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17972 13410 18000 15014
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14618 18184 14894
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18248 14482 18276 15150
rect 18432 15026 18460 16050
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18328 14408 18380 14414
rect 18328 14350 18380 14356
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17880 13382 18000 13410
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17236 12646 17264 13262
rect 17880 12866 17908 13382
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17972 12986 18000 13194
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17880 12838 18000 12866
rect 18156 12850 18184 13670
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12306 17264 12582
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17972 11694 18000 12838
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18340 12322 18368 14350
rect 18064 12294 18368 12322
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11286 17356 11494
rect 17420 11354 17448 11630
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17604 11370 17632 11562
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17512 11342 17632 11370
rect 17316 11280 17368 11286
rect 17316 11222 17368 11228
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9738 17264 9862
rect 17144 9710 17356 9738
rect 17144 9654 17172 9710
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 17040 9512 17092 9518
rect 16776 9438 16988 9466
rect 17040 9454 17092 9460
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 4554 16620 8978
rect 16684 8650 16712 9046
rect 16776 8974 16804 9438
rect 16960 9382 16988 9438
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16868 8974 16896 9318
rect 17052 9058 17080 9454
rect 17328 9110 17356 9710
rect 17316 9104 17368 9110
rect 17052 9042 17172 9058
rect 17316 9046 17368 9052
rect 17052 9036 17184 9042
rect 17052 9030 17132 9036
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16684 8634 16896 8650
rect 16684 8628 16908 8634
rect 16684 8622 16856 8628
rect 16856 8570 16908 8576
rect 16764 8560 16816 8566
rect 16684 8508 16764 8514
rect 16684 8502 16816 8508
rect 16684 8486 16804 8502
rect 16948 8492 17000 8498
rect 16684 8430 16712 8486
rect 16948 8434 17000 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16868 8090 16896 8366
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 6798 16712 7822
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16868 6934 16896 7482
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16960 6662 16988 8434
rect 17052 8430 17080 9030
rect 17132 8978 17184 8984
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 8430 17172 8502
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17236 8022 17264 8910
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7410 17172 7822
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17328 7546 17356 7754
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16592 3670 16620 4490
rect 16684 3942 16712 6598
rect 17328 6458 17356 6734
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16776 4826 16804 5170
rect 16764 4820 16816 4826
rect 16764 4762 16816 4768
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16408 2746 16528 2774
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16408 1834 16436 2746
rect 16396 1828 16448 1834
rect 16396 1770 16448 1776
rect 16776 800 16804 2790
rect 17144 2446 17172 3402
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17328 3126 17356 3334
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17236 800 17264 2790
rect 17328 2446 17356 3062
rect 17512 3058 17540 11342
rect 17696 10742 17724 11630
rect 18064 11218 18092 12294
rect 18432 12238 18460 14962
rect 18524 13462 18552 15438
rect 18616 15434 18644 15506
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18616 14414 18644 15370
rect 18708 15026 18736 16050
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18800 15638 18828 15982
rect 18984 15910 19012 15982
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18984 15502 19012 15846
rect 19076 15706 19104 16050
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 15706 19196 15914
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19076 15570 19104 15642
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 19260 15434 19288 15846
rect 20260 15632 20312 15638
rect 20258 15600 20260 15609
rect 20312 15600 20314 15609
rect 20258 15535 20314 15544
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 20364 15366 20392 15846
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 20916 15026 20944 16118
rect 21640 15088 21692 15094
rect 21638 15056 21640 15065
rect 21692 15056 21694 15065
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 20904 15020 20956 15026
rect 21638 14991 21694 15000
rect 20904 14962 20956 14968
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18800 14822 18828 14894
rect 18788 14816 18840 14822
rect 20916 14793 20944 14962
rect 21640 14952 21692 14958
rect 21638 14920 21640 14929
rect 21692 14920 21694 14929
rect 21638 14855 21694 14864
rect 21640 14816 21692 14822
rect 18788 14758 18840 14764
rect 20902 14784 20958 14793
rect 21744 14804 21772 17031
rect 21836 15162 21864 22066
rect 22112 21894 22140 22986
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23032 22234 23060 22578
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23400 22166 23428 22374
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22388 21622 22416 21966
rect 22376 21616 22428 21622
rect 22296 21564 22376 21570
rect 22296 21558 22428 21564
rect 22296 21542 22416 21558
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 22020 20534 22048 20810
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 19922 22232 20402
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 18970 22140 19314
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22020 17762 22048 18226
rect 22204 18086 22232 18770
rect 22296 18154 22324 21542
rect 22376 21412 22428 21418
rect 22376 21354 22428 21360
rect 22388 20806 22416 21354
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 20602 22416 20742
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22480 20466 22508 21966
rect 23020 21888 23072 21894
rect 23124 21876 23152 21966
rect 23400 21962 23428 22102
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23296 21888 23348 21894
rect 23124 21848 23296 21876
rect 23020 21830 23072 21836
rect 23296 21830 23348 21836
rect 23032 20874 23060 21830
rect 24688 21486 24716 23054
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24780 21690 24808 22646
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 23032 19990 23060 20810
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23400 20330 23428 20742
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 24122 20088 24178 20097
rect 24122 20023 24124 20032
rect 24176 20023 24178 20032
rect 24124 19994 24176 20000
rect 23020 19984 23072 19990
rect 23020 19926 23072 19932
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22388 18970 22416 19722
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22388 18766 22416 18906
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22376 18352 22428 18358
rect 22376 18294 22428 18300
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22020 17734 22140 17762
rect 21916 17604 21968 17610
rect 21916 17546 21968 17552
rect 21928 17134 21956 17546
rect 22112 17134 22140 17734
rect 22388 17542 22416 18294
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22388 17338 22416 17478
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 22112 16454 22140 16662
rect 22204 16658 22232 17274
rect 22282 17232 22338 17241
rect 22282 17167 22284 17176
rect 22336 17167 22338 17176
rect 22284 17138 22336 17144
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15434 21956 16050
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22020 15502 22048 15846
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 22112 15348 22140 16390
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15502 22232 15846
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22112 15320 22232 15348
rect 21824 15156 21876 15162
rect 22100 15156 22152 15162
rect 21876 15116 22100 15144
rect 21824 15098 21876 15104
rect 22100 15098 22152 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21692 14776 21772 14804
rect 21640 14758 21692 14764
rect 20902 14719 20958 14728
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18524 12986 18552 13398
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18156 11762 18184 12174
rect 18616 11762 18644 14350
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 20272 13938 20300 14282
rect 21376 14074 21404 14350
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12986 18736 13126
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18052 11212 18104 11218
rect 18052 11154 18104 11160
rect 17684 10736 17736 10742
rect 17736 10696 17908 10724
rect 17684 10678 17736 10684
rect 17880 9568 17908 10696
rect 18064 10266 18092 11154
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17604 9540 17908 9568
rect 17604 8430 17632 9540
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17696 7954 17724 9386
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9042 17816 9318
rect 17880 9178 17908 9540
rect 18064 9518 18092 10202
rect 18248 10062 18276 11630
rect 18616 11218 18644 11698
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18236 9716 18288 9722
rect 18340 9704 18368 11154
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18432 10713 18460 11086
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 19168 10538 19196 12786
rect 19260 12782 19288 13670
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19444 12918 19472 13262
rect 19982 13152 20038 13161
rect 19574 13084 19882 13104
rect 19982 13087 20038 13096
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19996 12918 20024 13087
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 20088 12434 20116 13262
rect 19996 12406 20116 12434
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11257 19472 12242
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19430 11248 19486 11257
rect 19352 11206 19430 11234
rect 19248 11144 19300 11150
rect 19352 11132 19380 11206
rect 19430 11183 19486 11192
rect 19300 11104 19380 11132
rect 19248 11086 19300 11092
rect 19524 11076 19576 11082
rect 19444 11036 19524 11064
rect 19338 10976 19394 10985
rect 19338 10911 19394 10920
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18288 9676 18368 9704
rect 18236 9658 18288 9664
rect 18248 9586 18276 9658
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18432 9518 18460 9862
rect 19352 9586 19380 10911
rect 19444 10742 19472 11036
rect 19524 11018 19576 11024
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10736 19484 10742
rect 19524 10736 19576 10742
rect 19432 10678 19484 10684
rect 19522 10704 19524 10713
rect 19576 10704 19578 10713
rect 19522 10639 19578 10648
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19536 10062 19564 10542
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18420 9512 18472 9518
rect 19352 9489 19380 9522
rect 18420 9454 18472 9460
rect 19338 9480 19394 9489
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17696 6798 17724 7346
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17788 5370 17816 7686
rect 17880 6662 17908 8910
rect 18432 7954 18460 9454
rect 19338 9415 19394 9424
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 19352 7886 19380 9415
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17788 4554 17816 5306
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19076 3942 19104 4082
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17696 800 17724 3334
rect 18524 2446 18552 3334
rect 18800 2774 18828 3470
rect 18984 3126 19012 3878
rect 19260 3398 19288 7414
rect 19352 5234 19380 7822
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19444 6322 19472 6938
rect 19904 6798 19932 7278
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19996 6390 20024 12406
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20088 9178 20116 9522
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19984 6384 20036 6390
rect 19890 6352 19946 6361
rect 19432 6316 19484 6322
rect 19984 6326 20036 6332
rect 19890 6287 19946 6296
rect 19432 6258 19484 6264
rect 19444 5642 19472 6258
rect 19904 5846 19932 6287
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5914 20024 6054
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19524 4752 19576 4758
rect 19524 4694 19576 4700
rect 19536 4554 19564 4694
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4146 19472 4422
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19996 3194 20024 5646
rect 20088 3194 20116 6666
rect 20180 6458 20208 13330
rect 20272 13326 20300 13874
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20824 12918 20852 13670
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20364 11286 20392 11834
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11354 20944 11698
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10742 20668 10950
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 9042 20668 9318
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20628 8900 20680 8906
rect 20628 8842 20680 8848
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20640 7410 20668 8842
rect 20732 8634 20760 8842
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20824 7546 20852 7754
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20260 6792 20312 6798
rect 20312 6740 20668 6746
rect 20260 6734 20668 6740
rect 20272 6730 20668 6734
rect 20272 6724 20680 6730
rect 20272 6718 20628 6724
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20272 6202 20300 6718
rect 20628 6666 20680 6672
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6322 20576 6598
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20180 6174 20300 6202
rect 20732 6186 20760 7278
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20720 6180 20772 6186
rect 20180 5710 20208 6174
rect 20720 6122 20772 6128
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20272 4622 20300 6054
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20640 5778 20668 5850
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20824 5370 20852 6190
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20444 4548 20496 4554
rect 20444 4490 20496 4496
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20180 3670 20208 4218
rect 20260 3936 20312 3942
rect 20258 3904 20260 3913
rect 20352 3936 20404 3942
rect 20312 3904 20314 3913
rect 20352 3878 20404 3884
rect 20258 3839 20314 3848
rect 20168 3664 20220 3670
rect 20168 3606 20220 3612
rect 20364 3602 20392 3878
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18708 2746 18828 2774
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18708 800 18736 2746
rect 19352 2650 19380 3130
rect 20272 3058 20300 3470
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 19076 2378 19104 2479
rect 19064 2372 19116 2378
rect 19064 2314 19116 2320
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19168 800 19196 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19720 870 19840 898
rect 19720 800 19748 870
rect 9048 734 9260 762
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 19812 762 19840 870
rect 19996 762 20024 2246
rect 20456 1902 20484 4490
rect 20548 3534 20576 5170
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20916 2514 20944 11290
rect 21192 10062 21220 12582
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11898 21312 12174
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21376 9110 21404 14010
rect 21468 14006 21496 14214
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21652 13705 21680 13738
rect 21638 13696 21694 13705
rect 21638 13631 21694 13640
rect 21744 13394 21772 14776
rect 21824 14816 21876 14822
rect 22112 14793 22140 14962
rect 21824 14758 21876 14764
rect 22098 14784 22154 14793
rect 21836 13734 21864 14758
rect 22098 14719 22154 14728
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21928 13546 21956 13874
rect 21836 13518 21956 13546
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21468 12986 21496 13262
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21468 12306 21496 12922
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21468 11642 21496 11698
rect 21640 11688 21692 11694
rect 21638 11656 21640 11665
rect 21692 11656 21694 11665
rect 21468 11614 21588 11642
rect 21560 11082 21588 11614
rect 21638 11591 21694 11600
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21376 8362 21404 8910
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21560 8090 21588 11018
rect 21744 8906 21772 13330
rect 21836 11762 21864 13518
rect 22112 13326 22140 14719
rect 22204 14346 22232 15320
rect 22282 15056 22338 15065
rect 22480 15026 22508 19858
rect 24412 19854 24440 21422
rect 25240 21146 25268 21490
rect 25228 21140 25280 21146
rect 25228 21082 25280 21088
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18834 22600 19110
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22572 18630 22600 18770
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22664 17202 22692 18702
rect 24412 18630 24440 19790
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24688 19514 24716 19722
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19514 25084 19654
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25148 18902 25176 19314
rect 25516 19242 25544 27338
rect 27068 25492 27120 25498
rect 27068 25434 27120 25440
rect 25780 23044 25832 23050
rect 25780 22986 25832 22992
rect 25792 22778 25820 22986
rect 26792 22976 26844 22982
rect 26792 22918 26844 22924
rect 26804 22778 26832 22918
rect 25780 22772 25832 22778
rect 25780 22714 25832 22720
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22030 26280 22578
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 25976 21146 26004 21286
rect 25964 21140 26016 21146
rect 25964 21082 26016 21088
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25792 20602 25820 20878
rect 26068 20806 26096 21286
rect 26252 20942 26280 21966
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26160 19718 26188 20402
rect 26240 19780 26292 19786
rect 26240 19722 26292 19728
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25412 18896 25464 18902
rect 25412 18838 25464 18844
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 17746 24440 18566
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 24400 17740 24452 17746
rect 24400 17682 24452 17688
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22664 15502 22692 17138
rect 23952 16114 23980 17682
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24688 17338 24716 17546
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 24688 16726 24716 17002
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24136 16182 24164 16526
rect 24124 16176 24176 16182
rect 24124 16118 24176 16124
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22282 14991 22338 15000
rect 22468 15020 22520 15026
rect 22296 14890 22324 14991
rect 22468 14962 22520 14968
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 23204 14476 23256 14482
rect 23204 14418 23256 14424
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12458 22140 12582
rect 21928 12442 22140 12458
rect 21916 12436 22140 12442
rect 21968 12430 22140 12436
rect 21916 12378 21968 12384
rect 21928 12347 21956 12378
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22112 12102 22140 12242
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22204 11914 22232 14282
rect 22836 13524 22888 13530
rect 22836 13466 22888 13472
rect 22848 13326 22876 13466
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22112 11886 22232 11914
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 22008 9512 22060 9518
rect 22006 9480 22008 9489
rect 22060 9480 22062 9489
rect 22006 9415 22062 9424
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 22112 8634 22140 11886
rect 22374 11656 22430 11665
rect 22374 11591 22430 11600
rect 22388 11354 22416 11591
rect 22572 11354 22600 12582
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22652 12164 22704 12170
rect 22652 12106 22704 12112
rect 22664 11801 22692 12106
rect 22756 11830 22784 12310
rect 22744 11824 22796 11830
rect 22650 11792 22706 11801
rect 22744 11766 22796 11772
rect 22650 11727 22706 11736
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22204 9058 22232 11222
rect 22296 11082 22324 11222
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22388 10810 22416 11290
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22388 9178 22416 9522
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22204 9030 22416 9058
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21178 7848 21234 7857
rect 21178 7783 21234 7792
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21008 6934 21036 7686
rect 20996 6928 21048 6934
rect 20994 6896 20996 6905
rect 21048 6896 21050 6905
rect 20994 6831 21050 6840
rect 21192 5574 21220 7783
rect 21560 7002 21588 8026
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21284 5370 21312 6598
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21468 5846 21496 6258
rect 21652 6118 21680 6938
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21744 5778 21772 8298
rect 22192 7812 22244 7818
rect 22192 7754 22244 7760
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7342 21864 7686
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21928 6866 21956 7142
rect 22204 6866 22232 7754
rect 22282 6896 22338 6905
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 22192 6860 22244 6866
rect 22282 6831 22338 6840
rect 22192 6802 22244 6808
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21836 5302 21864 6054
rect 21928 5710 21956 6802
rect 22296 6798 22324 6831
rect 22388 6798 22416 9030
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22756 7410 22784 7822
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22480 6730 22508 7346
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22848 6322 22876 13262
rect 22940 13190 22968 14350
rect 23032 14074 23060 14350
rect 23216 14074 23244 14418
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22940 12238 22968 13126
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 12102 23060 12174
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23308 11880 23336 14962
rect 23952 13938 23980 16050
rect 24596 15706 24624 16050
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 24136 12374 24164 15642
rect 24872 15570 24900 16526
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24964 15502 24992 16186
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25056 14482 25084 17070
rect 25148 16590 25176 18634
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 17134 25268 17478
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25332 16454 25360 17070
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 25424 15502 25452 18838
rect 26160 18698 26188 19654
rect 26252 19446 26280 19722
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26252 18748 26280 19382
rect 26436 19174 26464 22646
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26252 18720 26556 18748
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 25686 17504 25742 17513
rect 25686 17439 25742 17448
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25516 17134 25544 17274
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25700 17066 25728 17439
rect 26252 17202 26280 17818
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26068 17105 26096 17138
rect 26054 17096 26110 17105
rect 25688 17060 25740 17066
rect 26054 17031 26110 17040
rect 25688 17002 25740 17008
rect 26068 16658 26096 17031
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26528 16590 26556 18720
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 24412 13190 24440 14010
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24412 12617 24440 12718
rect 24398 12608 24454 12617
rect 24398 12543 24454 12552
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 22940 11852 23336 11880
rect 22940 7206 22968 11852
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23032 11150 23060 11698
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23124 11354 23152 11494
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23216 11286 23244 11562
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 23308 11014 23336 11562
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23400 10810 23428 11086
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23492 9518 23520 9549
rect 23480 9512 23532 9518
rect 23478 9480 23480 9489
rect 23532 9480 23534 9489
rect 23478 9415 23534 9424
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 8906 23152 9318
rect 23112 8900 23164 8906
rect 23112 8842 23164 8848
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23216 8634 23244 8842
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23492 7342 23520 9415
rect 23584 9110 23612 12106
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23584 8498 23612 9046
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 22928 7200 22980 7206
rect 22928 7142 22980 7148
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 22112 5846 22140 6190
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22204 5914 22232 6122
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 22100 5840 22152 5846
rect 22100 5782 22152 5788
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21824 5296 21876 5302
rect 21824 5238 21876 5244
rect 22296 4690 22324 6190
rect 22480 6118 22508 6190
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 23492 5778 23520 7278
rect 23480 5772 23532 5778
rect 23480 5714 23532 5720
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 23294 5128 23350 5137
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22006 4040 22062 4049
rect 22112 4010 22140 4422
rect 22480 4078 22508 5102
rect 23294 5063 23350 5072
rect 23308 4690 23336 5063
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22376 4072 22428 4078
rect 22190 4040 22246 4049
rect 22006 3975 22062 3984
rect 22100 4004 22152 4010
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 21100 3194 21128 3402
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21836 3058 21864 3606
rect 22020 3126 22048 3975
rect 22376 4014 22428 4020
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22190 3975 22192 3984
rect 22100 3946 22152 3952
rect 22244 3975 22246 3984
rect 22192 3946 22244 3952
rect 22098 3768 22154 3777
rect 22098 3703 22154 3712
rect 22112 3670 22140 3703
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22008 3120 22060 3126
rect 22008 3062 22060 3068
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20180 870 20300 898
rect 20180 800 20208 870
rect 19812 734 20024 762
rect 20166 0 20222 800
rect 20272 762 20300 870
rect 20548 762 20576 2246
rect 21100 800 21128 2994
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21652 800 21680 2790
rect 22020 2038 22048 3062
rect 22204 2650 22232 3606
rect 22388 3194 22416 4014
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22480 3074 22508 4014
rect 22664 3534 22692 4558
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23032 3670 23060 4014
rect 23308 3670 23336 4082
rect 23020 3664 23072 3670
rect 22926 3632 22982 3641
rect 23020 3606 23072 3612
rect 23296 3664 23348 3670
rect 23296 3606 23348 3612
rect 22926 3567 22982 3576
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22388 3046 22508 3074
rect 22664 3058 22692 3470
rect 22652 3052 22704 3058
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22100 2576 22152 2582
rect 22100 2518 22152 2524
rect 22008 2032 22060 2038
rect 22008 1974 22060 1980
rect 22112 800 22140 2518
rect 22388 2514 22416 3046
rect 22652 2994 22704 3000
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22480 2650 22508 2926
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22664 1442 22692 2858
rect 22756 2666 22784 3470
rect 22940 3466 22968 3567
rect 23032 3534 23060 3606
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 22940 3058 22968 3402
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 3126 23060 3334
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23492 3058 23520 3470
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 22756 2650 22876 2666
rect 22756 2644 22888 2650
rect 22756 2638 22836 2644
rect 22756 1494 22784 2638
rect 22836 2586 22888 2592
rect 22940 2446 22968 2790
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23216 2106 23244 2382
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 22572 1414 22692 1442
rect 22744 1488 22796 1494
rect 22744 1430 22796 1436
rect 22572 800 22600 1414
rect 23584 800 23612 4082
rect 23676 4010 23704 10950
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23768 8498 23796 8978
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23768 7478 23796 8230
rect 23860 7750 23888 8366
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 24412 6390 24440 12543
rect 24504 11150 24532 14010
rect 25884 13802 25912 14350
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25688 13728 25740 13734
rect 25688 13670 25740 13676
rect 25700 13530 25728 13670
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24688 12714 24716 13262
rect 24872 12986 24900 13262
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24124 5772 24176 5778
rect 24124 5714 24176 5720
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 24136 3058 24164 5714
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24228 4826 24256 5170
rect 24504 5166 24532 11086
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24596 8566 24624 8910
rect 24584 8560 24636 8566
rect 24584 8502 24636 8508
rect 24596 5681 24624 8502
rect 24582 5672 24638 5681
rect 24582 5607 24638 5616
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 23768 2854 23796 2994
rect 23756 2848 23808 2854
rect 23756 2790 23808 2796
rect 24320 2378 24348 4490
rect 24504 4282 24532 4558
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24412 3602 24440 4082
rect 24504 3670 24532 4218
rect 24688 4185 24716 12650
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25332 11898 25360 12174
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25240 11354 25268 11766
rect 25332 11762 25360 11834
rect 25608 11830 25636 12038
rect 25976 11898 26004 14554
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26068 12850 26096 13670
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 26068 12434 26096 12786
rect 26160 12646 26188 16526
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26344 15434 26372 15914
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26436 15706 26464 15846
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26528 15434 26556 16526
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26620 15570 26648 15642
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26516 15428 26568 15434
rect 26516 15370 26568 15376
rect 26528 14482 26556 15370
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26620 14414 26648 14894
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26148 12640 26200 12646
rect 26148 12582 26200 12588
rect 26068 12406 26188 12434
rect 26160 12238 26188 12406
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25964 11892 26016 11898
rect 25964 11834 26016 11840
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 25596 11824 25648 11830
rect 25596 11766 25648 11772
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25504 11280 25556 11286
rect 25424 11228 25504 11234
rect 25424 11222 25556 11228
rect 25424 11206 25544 11222
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 25148 7206 25176 7754
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 7002 25176 7142
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24872 5370 24900 5578
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 24780 4570 24808 5034
rect 24860 4616 24912 4622
rect 24780 4564 24860 4570
rect 24780 4558 24912 4564
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 24780 4542 24900 4558
rect 24674 4176 24730 4185
rect 24674 4111 24730 4120
rect 24492 3664 24544 3670
rect 24780 3618 24808 4542
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24492 3606 24544 3612
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24596 3590 24808 3618
rect 24492 3528 24544 3534
rect 24596 3516 24624 3590
rect 24872 3534 24900 4150
rect 24544 3488 24624 3516
rect 24860 3528 24912 3534
rect 24492 3470 24544 3476
rect 24860 3470 24912 3476
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24872 2446 24900 3130
rect 25148 2854 25176 4558
rect 25424 3777 25452 11206
rect 25596 6112 25648 6118
rect 25596 6054 25648 6060
rect 25608 5234 25636 6054
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25504 4140 25556 4146
rect 25608 4128 25636 5170
rect 25556 4100 25636 4128
rect 25504 4082 25556 4088
rect 25410 3768 25466 3777
rect 25410 3703 25466 3712
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 25424 3126 25452 3334
rect 25608 3194 25636 3470
rect 25700 3194 25728 11698
rect 25792 11558 25820 11698
rect 26068 11626 26096 11834
rect 26160 11762 26188 12174
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26056 11620 26108 11626
rect 26056 11562 26108 11568
rect 25780 11552 25832 11558
rect 25780 11494 25832 11500
rect 25792 11082 25820 11494
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 25872 9920 25924 9926
rect 25872 9862 25924 9868
rect 25884 9654 25912 9862
rect 25872 9648 25924 9654
rect 25872 9590 25924 9596
rect 26068 9042 26096 11562
rect 26160 11286 26188 11698
rect 26148 11280 26200 11286
rect 26148 11222 26200 11228
rect 26344 11150 26372 13806
rect 26620 13326 26648 14350
rect 26804 13462 26832 20810
rect 27080 19174 27108 25434
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 28000 22778 28028 23054
rect 28448 22976 28500 22982
rect 28448 22918 28500 22924
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 28460 22710 28488 22918
rect 28448 22704 28500 22710
rect 28448 22646 28500 22652
rect 31220 22642 31248 23054
rect 31484 23044 31536 23050
rect 31484 22986 31536 22992
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 27632 22234 27660 22578
rect 27896 22568 27948 22574
rect 27896 22510 27948 22516
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27264 20874 27292 21286
rect 27620 20936 27672 20942
rect 27620 20878 27672 20884
rect 27252 20868 27304 20874
rect 27252 20810 27304 20816
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27172 20058 27200 20402
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27172 19446 27200 19722
rect 27356 19514 27384 20402
rect 27540 19786 27568 20742
rect 27632 20602 27660 20878
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27724 20398 27752 20538
rect 27908 20398 27936 22510
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28460 22001 28488 22170
rect 30208 22166 30236 22374
rect 28816 22160 28868 22166
rect 28816 22102 28868 22108
rect 28908 22160 28960 22166
rect 28908 22102 28960 22108
rect 30196 22160 30248 22166
rect 30196 22102 30248 22108
rect 28446 21992 28502 22001
rect 28446 21927 28502 21936
rect 28828 21554 28856 22102
rect 28920 21690 28948 22102
rect 30208 22030 30236 22102
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 28908 21684 28960 21690
rect 28908 21626 28960 21632
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28828 21350 28856 21490
rect 28264 21344 28316 21350
rect 28264 21286 28316 21292
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28276 21010 28304 21286
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 28264 21004 28316 21010
rect 28264 20946 28316 20952
rect 28092 20806 28120 20946
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 28000 20534 28028 20742
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27896 20392 27948 20398
rect 27896 20334 27948 20340
rect 27528 19780 27580 19786
rect 27528 19722 27580 19728
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27160 19440 27212 19446
rect 27160 19382 27212 19388
rect 27540 19360 27568 19722
rect 27540 19332 27660 19360
rect 27068 19168 27120 19174
rect 27068 19110 27120 19116
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 27080 18290 27108 18566
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27080 17762 27108 18226
rect 27172 17882 27200 18226
rect 27160 17876 27212 17882
rect 27160 17818 27212 17824
rect 27080 17734 27292 17762
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 27080 17338 27108 17614
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26436 11558 26464 12174
rect 26528 12102 26556 13126
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26896 10198 26924 17138
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27172 15162 27200 15370
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27080 14278 27108 14962
rect 27264 14414 27292 17734
rect 27436 17740 27488 17746
rect 27436 17682 27488 17688
rect 27448 17202 27476 17682
rect 27526 17232 27582 17241
rect 27436 17196 27488 17202
rect 27526 17167 27528 17176
rect 27436 17138 27488 17144
rect 27580 17167 27582 17176
rect 27528 17138 27580 17144
rect 27448 16726 27476 17138
rect 27436 16720 27488 16726
rect 27436 16662 27488 16668
rect 27632 15026 27660 19332
rect 27908 18630 27936 20334
rect 28828 19854 28856 21286
rect 28906 20088 28962 20097
rect 28906 20023 28962 20032
rect 28920 19990 28948 20023
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28724 19440 28776 19446
rect 28724 19382 28776 19388
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 28000 15978 28028 19314
rect 28540 19304 28592 19310
rect 28540 19246 28592 19252
rect 27988 15972 28040 15978
rect 27988 15914 28040 15920
rect 27436 15020 27488 15026
rect 27436 14962 27488 14968
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27448 14618 27476 14962
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 27908 14618 27936 14758
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27264 13870 27292 14350
rect 28000 14006 28028 15914
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28276 15026 28304 15302
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28170 14920 28226 14929
rect 28170 14855 28226 14864
rect 28184 14822 28212 14855
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28092 14414 28120 14758
rect 28264 14544 28316 14550
rect 28264 14486 28316 14492
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28276 14278 28304 14486
rect 28264 14272 28316 14278
rect 28264 14214 28316 14220
rect 27988 14000 28040 14006
rect 27988 13942 28040 13948
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27908 13258 27936 13874
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 27896 13252 27948 13258
rect 27896 13194 27948 13200
rect 28000 12918 28028 13670
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28184 13161 28212 13194
rect 28170 13152 28226 13161
rect 28170 13087 28226 13096
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 28276 12850 28304 14214
rect 28356 13184 28408 13190
rect 28356 13126 28408 13132
rect 28368 12918 28396 13126
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27252 12164 27304 12170
rect 27252 12106 27304 12112
rect 26884 10192 26936 10198
rect 26884 10134 26936 10140
rect 26332 10056 26384 10062
rect 26332 9998 26384 10004
rect 26240 9444 26292 9450
rect 26240 9386 26292 9392
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 26252 8974 26280 9386
rect 26344 9178 26372 9998
rect 27068 9920 27120 9926
rect 27068 9862 27120 9868
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 7478 26740 7686
rect 26700 7472 26752 7478
rect 26700 7414 26752 7420
rect 26804 7342 26832 9454
rect 26896 9042 26924 9522
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26884 7880 26936 7886
rect 26882 7848 26884 7857
rect 26936 7848 26938 7857
rect 26882 7783 26938 7792
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25792 5234 25820 6394
rect 26068 6322 26096 6802
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26252 6322 26280 6598
rect 26804 6322 26832 7278
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 26792 6316 26844 6322
rect 26792 6258 26844 6264
rect 25884 6202 25912 6258
rect 25884 6174 26188 6202
rect 26160 6118 26188 6174
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26804 5710 26832 6258
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 26332 5636 26384 5642
rect 26332 5578 26384 5584
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25792 4282 25820 5170
rect 25884 5166 25912 5510
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25884 4554 25912 5102
rect 25872 4548 25924 4554
rect 25872 4490 25924 4496
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 25872 4140 25924 4146
rect 25792 4100 25872 4128
rect 25792 3466 25820 4100
rect 25976 4128 26004 5170
rect 26068 4758 26096 5510
rect 26344 5370 26372 5578
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 26160 4622 26188 5170
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 25924 4100 26004 4128
rect 25872 4082 25924 4088
rect 26896 3942 26924 7783
rect 27080 7750 27108 9862
rect 27160 8288 27212 8294
rect 27160 8230 27212 8236
rect 27172 7886 27200 8230
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27068 7744 27120 7750
rect 27068 7686 27120 7692
rect 26974 5672 27030 5681
rect 26974 5607 26976 5616
rect 27028 5607 27030 5616
rect 26976 5578 27028 5584
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26974 3904 27030 3913
rect 25872 3664 25924 3670
rect 25872 3606 25924 3612
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 25412 3120 25464 3126
rect 25412 3062 25464 3068
rect 25884 2854 25912 3606
rect 25976 3398 26004 3878
rect 26436 3534 26464 3878
rect 26974 3839 27030 3848
rect 26988 3670 27016 3839
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 27264 3194 27292 12106
rect 27448 11762 27476 12582
rect 28092 12220 28120 12786
rect 28172 12232 28224 12238
rect 28092 12192 28172 12220
rect 28092 11830 28120 12192
rect 28172 12174 28224 12180
rect 28080 11824 28132 11830
rect 28080 11766 28132 11772
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27356 10810 27384 11698
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27356 9450 27384 10746
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27540 7954 27568 8434
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27632 5846 27660 10610
rect 28172 9512 28224 9518
rect 28172 9454 28224 9460
rect 28184 8974 28212 9454
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 27804 8560 27856 8566
rect 27804 8502 27856 8508
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 27816 7954 27844 8502
rect 28080 8424 28132 8430
rect 28080 8366 28132 8372
rect 28092 8090 28120 8366
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27816 7750 27844 7890
rect 28184 7886 28212 8502
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 27712 7472 27764 7478
rect 27712 7414 27764 7420
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27632 5234 27660 5782
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27724 4486 27752 7414
rect 27816 7188 27844 7686
rect 28184 7410 28212 7686
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 27988 7200 28040 7206
rect 27816 7160 27988 7188
rect 27816 6361 27844 7160
rect 27988 7142 28040 7148
rect 27802 6352 27858 6361
rect 27802 6287 27858 6296
rect 27988 4548 28040 4554
rect 27988 4490 28040 4496
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 28000 3641 28028 4490
rect 27986 3632 28042 3641
rect 27986 3567 28042 3576
rect 27252 3188 27304 3194
rect 27252 3130 27304 3136
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 27436 3052 27488 3058
rect 27436 2994 27488 3000
rect 25136 2848 25188 2854
rect 25136 2790 25188 2796
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25608 2650 25636 2790
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24032 2304 24084 2310
rect 24676 2304 24728 2310
rect 24032 2246 24084 2252
rect 24596 2264 24676 2292
rect 24044 800 24072 2246
rect 24596 800 24624 2264
rect 24676 2246 24728 2252
rect 25056 800 25084 2518
rect 25976 800 26004 2994
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26528 800 26556 2246
rect 26896 2106 26924 2382
rect 26884 2100 26936 2106
rect 26884 2042 26936 2048
rect 27448 800 27476 2994
rect 28276 2446 28304 12786
rect 28460 11014 28488 12786
rect 28552 11801 28580 19246
rect 28736 18970 28764 19382
rect 28814 19272 28870 19281
rect 28814 19207 28870 19216
rect 28828 18970 28856 19207
rect 28906 19000 28962 19009
rect 28724 18964 28776 18970
rect 28724 18906 28776 18912
rect 28816 18964 28868 18970
rect 29012 18970 29040 19858
rect 29104 19718 29132 21966
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29196 21554 29224 21898
rect 30576 21690 30604 21966
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 31114 21584 31170 21593
rect 29184 21548 29236 21554
rect 31114 21519 31116 21528
rect 29184 21490 29236 21496
rect 31168 21519 31170 21528
rect 31116 21490 31168 21496
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29564 19854 29592 20198
rect 31220 19922 31248 22578
rect 31312 21418 31340 22578
rect 31496 22234 31524 22986
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32232 22710 32260 22918
rect 32220 22704 32272 22710
rect 32220 22646 32272 22652
rect 32404 22704 32456 22710
rect 32404 22646 32456 22652
rect 31760 22500 31812 22506
rect 31760 22442 31812 22448
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31392 22024 31444 22030
rect 31392 21966 31444 21972
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 29736 19916 29788 19922
rect 29736 19858 29788 19864
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29748 19718 29776 19858
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 29182 19272 29238 19281
rect 29182 19207 29238 19216
rect 28906 18935 28962 18944
rect 29000 18964 29052 18970
rect 28816 18906 28868 18912
rect 28920 18902 28948 18935
rect 29000 18906 29052 18912
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28644 18222 28672 18634
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 29012 17882 29040 18906
rect 29196 18766 29224 19207
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 18290 29224 18702
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28644 12646 28672 16050
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28816 14340 28868 14346
rect 28816 14282 28868 14288
rect 28736 13938 28764 14282
rect 28828 14074 28856 14282
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 28736 13326 28764 13874
rect 28814 13696 28870 13705
rect 28814 13631 28870 13640
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28538 11792 28594 11801
rect 28538 11727 28594 11736
rect 28552 11694 28580 11727
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 28736 11626 28764 12786
rect 28828 12714 28856 13631
rect 28920 13190 28948 17206
rect 29380 16726 29408 19110
rect 29472 18630 29500 19314
rect 29656 19281 29684 19314
rect 29642 19272 29698 19281
rect 29642 19207 29698 19216
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 18766 30052 19110
rect 30116 18834 30144 19654
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30208 18970 30236 19314
rect 30576 19310 30604 19790
rect 30760 19514 30788 19790
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30484 18970 30512 19246
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30104 18828 30156 18834
rect 30104 18770 30156 18776
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 29460 18624 29512 18630
rect 29460 18566 29512 18572
rect 29472 18290 29500 18566
rect 29564 18329 29592 18634
rect 29550 18320 29606 18329
rect 29460 18284 29512 18290
rect 29550 18255 29606 18264
rect 30380 18284 30432 18290
rect 29460 18226 29512 18232
rect 30380 18226 30432 18232
rect 30392 18154 30420 18226
rect 30288 18148 30340 18154
rect 30288 18090 30340 18096
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 29552 18080 29604 18086
rect 29552 18022 29604 18028
rect 29564 17678 29592 18022
rect 30300 17882 30328 18090
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 29552 17672 29604 17678
rect 29552 17614 29604 17620
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29368 16720 29420 16726
rect 29368 16662 29420 16668
rect 29840 16522 29868 17138
rect 30300 17134 30328 17274
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 29552 16516 29604 16522
rect 29552 16458 29604 16464
rect 29828 16516 29880 16522
rect 29828 16458 29880 16464
rect 29000 16448 29052 16454
rect 29000 16390 29052 16396
rect 29012 16114 29040 16390
rect 29380 16114 29408 16458
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29288 13870 29316 15982
rect 29564 15706 29592 16458
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29012 13394 29040 13738
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 29368 13320 29420 13326
rect 29368 13262 29420 13268
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 29276 13184 29328 13190
rect 29276 13126 29328 13132
rect 29288 12986 29316 13126
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29380 12850 29408 13262
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28954 12640 29006 12646
rect 28814 12608 28870 12617
rect 28870 12588 28954 12594
rect 28870 12582 29006 12588
rect 28870 12566 28994 12582
rect 28814 12543 28870 12552
rect 28724 11620 28776 11626
rect 28724 11562 28776 11568
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28736 7970 28764 8026
rect 28644 7942 28764 7970
rect 28644 7886 28672 7942
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28644 7478 28672 7822
rect 28632 7472 28684 7478
rect 28632 7414 28684 7420
rect 28920 2650 28948 10950
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29564 9382 29592 9522
rect 29552 9376 29604 9382
rect 29552 9318 29604 9324
rect 29564 7818 29592 9318
rect 29552 7812 29604 7818
rect 29552 7754 29604 7760
rect 29552 6792 29604 6798
rect 29552 6734 29604 6740
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29104 5778 29132 6258
rect 29564 5778 29592 6734
rect 29736 6316 29788 6322
rect 29736 6258 29788 6264
rect 29748 6225 29776 6258
rect 29734 6216 29790 6225
rect 29734 6151 29790 6160
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 29552 5772 29604 5778
rect 29552 5714 29604 5720
rect 29000 4752 29052 4758
rect 29000 4694 29052 4700
rect 29012 4146 29040 4694
rect 29104 4214 29132 5714
rect 29656 5710 29684 6054
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29104 3058 29132 4150
rect 29564 4078 29592 4558
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29564 3942 29592 4014
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 29564 2446 29592 3878
rect 29840 3097 29868 16458
rect 30288 15904 30340 15910
rect 30208 15864 30288 15892
rect 30208 15502 30236 15864
rect 30288 15846 30340 15852
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30300 14090 30328 15438
rect 30392 15434 30420 16526
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30392 15162 30420 15370
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30392 14482 30420 15098
rect 30484 15026 30512 16118
rect 30576 15502 30604 17614
rect 30564 15496 30616 15502
rect 30668 15484 30696 19314
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 30838 18456 30894 18465
rect 30838 18391 30894 18400
rect 30852 18358 30880 18391
rect 30840 18352 30892 18358
rect 30840 18294 30892 18300
rect 30944 18290 30972 18702
rect 31128 18290 31156 19314
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 30944 17202 30972 18226
rect 31220 17746 31248 18294
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 15638 30788 16390
rect 30944 15910 30972 16526
rect 31128 16250 31156 17138
rect 31208 16516 31260 16522
rect 31208 16458 31260 16464
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31128 16114 31156 16186
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 30932 15904 30984 15910
rect 30932 15846 30984 15852
rect 30748 15632 30800 15638
rect 30748 15574 30800 15580
rect 30668 15456 30788 15484
rect 30564 15438 30616 15444
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30380 14476 30432 14482
rect 30380 14418 30432 14424
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30116 14062 30328 14090
rect 30116 13530 30144 14062
rect 30392 14006 30420 14214
rect 30380 14000 30432 14006
rect 30286 13968 30342 13977
rect 30380 13942 30432 13948
rect 30286 13903 30288 13912
rect 30340 13903 30342 13912
rect 30288 13874 30340 13880
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 29932 11830 29960 13466
rect 30104 12912 30156 12918
rect 30104 12854 30156 12860
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 30012 8968 30064 8974
rect 30012 8910 30064 8916
rect 30024 8430 30052 8910
rect 30012 8424 30064 8430
rect 30012 8366 30064 8372
rect 30010 6488 30066 6497
rect 30010 6423 30012 6432
rect 30064 6423 30066 6432
rect 30012 6394 30064 6400
rect 29826 3088 29882 3097
rect 29826 3023 29882 3032
rect 30116 2650 30144 12854
rect 30208 12306 30236 13806
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30208 11218 30236 12242
rect 30484 11898 30512 14962
rect 30656 14068 30708 14074
rect 30656 14010 30708 14016
rect 30668 13326 30696 14010
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30760 12434 30788 15456
rect 31220 15366 31248 16458
rect 31312 15434 31340 17138
rect 31300 15428 31352 15434
rect 31300 15370 31352 15376
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 31208 15360 31260 15366
rect 31208 15302 31260 15308
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30944 14958 30972 15030
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30852 13530 30880 14350
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 30944 13326 30972 14894
rect 31036 14482 31064 15302
rect 31404 15178 31432 21966
rect 31484 21956 31536 21962
rect 31484 21898 31536 21904
rect 31496 21842 31524 21898
rect 31772 21842 31800 22442
rect 31944 22432 31996 22438
rect 31944 22374 31996 22380
rect 31956 22030 31984 22374
rect 32036 22160 32088 22166
rect 32036 22102 32088 22108
rect 31944 22024 31996 22030
rect 31944 21966 31996 21972
rect 31496 21814 31800 21842
rect 31852 21888 31904 21894
rect 31852 21830 31904 21836
rect 31496 21690 31524 21814
rect 31484 21684 31536 21690
rect 31484 21626 31536 21632
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31588 20942 31616 21626
rect 31864 21350 31892 21830
rect 32048 21622 32076 22102
rect 32036 21616 32088 21622
rect 32232 21593 32260 22646
rect 32036 21558 32088 21564
rect 32218 21584 32274 21593
rect 32218 21519 32274 21528
rect 32416 21486 32444 22646
rect 32404 21480 32456 21486
rect 32404 21422 32456 21428
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 31588 19310 31616 20878
rect 32048 19378 32168 19394
rect 32036 19372 32168 19378
rect 32088 19366 32168 19372
rect 32036 19314 32088 19320
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31944 19236 31996 19242
rect 31944 19178 31996 19184
rect 32036 19236 32088 19242
rect 32036 19178 32088 19184
rect 31852 18828 31904 18834
rect 31852 18770 31904 18776
rect 31576 18352 31628 18358
rect 31576 18294 31628 18300
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31496 17882 31524 18022
rect 31484 17876 31536 17882
rect 31484 17818 31536 17824
rect 31484 15428 31536 15434
rect 31484 15370 31536 15376
rect 31312 15150 31432 15178
rect 31208 14612 31260 14618
rect 31208 14554 31260 14560
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 31036 14278 31064 14418
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31128 12646 31156 14350
rect 31116 12640 31168 12646
rect 31116 12582 31168 12588
rect 30760 12406 31064 12434
rect 30472 11892 30524 11898
rect 30472 11834 30524 11840
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30208 9382 30236 10542
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 30208 8294 30236 9318
rect 30300 8362 30328 11494
rect 30668 11354 30696 11766
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30932 8900 30984 8906
rect 30932 8842 30984 8848
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30300 8022 30328 8298
rect 30288 8016 30340 8022
rect 30288 7958 30340 7964
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30484 6322 30512 7822
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30484 4622 30512 4966
rect 30668 4826 30696 6326
rect 30656 4820 30708 4826
rect 30656 4762 30708 4768
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30196 4548 30248 4554
rect 30196 4490 30248 4496
rect 30208 3942 30236 4490
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30300 2990 30328 4082
rect 30852 3058 30880 8774
rect 30944 8634 30972 8842
rect 31036 8634 31064 12406
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 30932 8628 30984 8634
rect 30932 8570 30984 8576
rect 31024 8628 31076 8634
rect 31024 8570 31076 8576
rect 31128 8498 31156 9318
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31220 8344 31248 14554
rect 31128 8316 31248 8344
rect 30932 7336 30984 7342
rect 30932 7278 30984 7284
rect 30944 6866 30972 7278
rect 30932 6860 30984 6866
rect 30932 6802 30984 6808
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 30932 6384 30984 6390
rect 30932 6326 30984 6332
rect 30944 5846 30972 6326
rect 31036 6322 31064 6734
rect 31128 6458 31156 8316
rect 31312 7970 31340 15150
rect 31390 14920 31446 14929
rect 31390 14855 31446 14864
rect 31404 14618 31432 14855
rect 31392 14612 31444 14618
rect 31392 14554 31444 14560
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31404 14074 31432 14350
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31220 7942 31340 7970
rect 31116 6452 31168 6458
rect 31116 6394 31168 6400
rect 31024 6316 31076 6322
rect 31024 6258 31076 6264
rect 30932 5840 30984 5846
rect 30932 5782 30984 5788
rect 30944 4554 30972 5782
rect 31116 4616 31168 4622
rect 31114 4584 31116 4593
rect 31168 4584 31170 4593
rect 30932 4548 30984 4554
rect 31114 4519 31170 4528
rect 30932 4490 30984 4496
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 30300 2854 30328 2926
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 30300 2514 30328 2790
rect 30852 2582 30880 2994
rect 30840 2576 30892 2582
rect 30840 2518 30892 2524
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 30944 2446 30972 4490
rect 31128 3534 31156 4519
rect 31220 3602 31248 7942
rect 31404 6662 31432 8230
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31300 4548 31352 4554
rect 31300 4490 31352 4496
rect 31312 4282 31340 4490
rect 31300 4276 31352 4282
rect 31300 4218 31352 4224
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31022 3224 31078 3233
rect 31022 3159 31024 3168
rect 31076 3159 31078 3168
rect 31024 3130 31076 3136
rect 31128 3058 31156 3334
rect 31220 3194 31248 3402
rect 31496 3210 31524 15370
rect 31588 11064 31616 18294
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31680 17134 31708 18226
rect 31864 17746 31892 18770
rect 31852 17740 31904 17746
rect 31852 17682 31904 17688
rect 31864 17270 31892 17682
rect 31852 17264 31904 17270
rect 31852 17206 31904 17212
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31852 16720 31904 16726
rect 31852 16662 31904 16668
rect 31760 14952 31812 14958
rect 31758 14920 31760 14929
rect 31812 14920 31814 14929
rect 31758 14855 31814 14864
rect 31668 14544 31720 14550
rect 31668 14486 31720 14492
rect 31680 14414 31708 14486
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31680 13190 31708 14350
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31760 12164 31812 12170
rect 31760 12106 31812 12112
rect 31588 11036 31708 11064
rect 31576 10532 31628 10538
rect 31576 10474 31628 10480
rect 31588 9926 31616 10474
rect 31576 9920 31628 9926
rect 31576 9862 31628 9868
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 31588 4486 31616 4558
rect 31680 4536 31708 11036
rect 31772 9518 31800 12106
rect 31864 10010 31892 16662
rect 31956 10130 31984 19178
rect 32048 18766 32076 19178
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 32048 17814 32076 18702
rect 32140 18222 32168 19366
rect 32220 19304 32272 19310
rect 32218 19272 32220 19281
rect 32272 19272 32274 19281
rect 32218 19207 32274 19216
rect 32232 18766 32260 19207
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32128 18216 32180 18222
rect 32128 18158 32180 18164
rect 32036 17808 32088 17814
rect 32036 17750 32088 17756
rect 32048 17202 32076 17750
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32140 16182 32168 18158
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32416 17218 32444 17614
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 32324 17190 32444 17218
rect 32128 16176 32180 16182
rect 32128 16118 32180 16124
rect 32232 15994 32260 17138
rect 32140 15978 32260 15994
rect 32128 15972 32260 15978
rect 32180 15966 32260 15972
rect 32128 15914 32180 15920
rect 32140 15502 32168 15914
rect 32128 15496 32180 15502
rect 32128 15438 32180 15444
rect 32324 14890 32352 17190
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32416 15094 32444 16050
rect 32404 15088 32456 15094
rect 32404 15030 32456 15036
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32416 14618 32444 15030
rect 32404 14612 32456 14618
rect 32404 14554 32456 14560
rect 32128 13932 32180 13938
rect 32128 13874 32180 13880
rect 32140 13462 32168 13874
rect 32128 13456 32180 13462
rect 32128 13398 32180 13404
rect 32140 13326 32168 13398
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 32140 12238 32168 13262
rect 32508 12442 32536 38898
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34612 23112 34664 23118
rect 34612 23054 34664 23060
rect 34624 22642 34652 23054
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33968 22636 34020 22642
rect 33968 22578 34020 22584
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 32600 21962 32628 22578
rect 32772 22432 32824 22438
rect 32772 22374 32824 22380
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32588 21956 32640 21962
rect 32588 21898 32640 21904
rect 32692 21554 32720 21966
rect 32680 21548 32732 21554
rect 32680 21490 32732 21496
rect 32588 21480 32640 21486
rect 32588 21422 32640 21428
rect 32600 21010 32628 21422
rect 32784 21010 32812 22374
rect 33152 22098 33180 22578
rect 33140 22092 33192 22098
rect 33980 22094 34008 22578
rect 34716 22234 34744 22578
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 36268 22432 36320 22438
rect 36268 22374 36320 22380
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 33980 22066 34284 22094
rect 33140 22034 33192 22040
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33600 22024 33652 22030
rect 33600 21966 33652 21972
rect 33428 21690 33456 21966
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 32862 21584 32918 21593
rect 32862 21519 32864 21528
rect 32916 21519 32918 21528
rect 32864 21490 32916 21496
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 32588 21004 32640 21010
rect 32588 20946 32640 20952
rect 32772 21004 32824 21010
rect 32772 20946 32824 20952
rect 32588 19712 32640 19718
rect 32588 19654 32640 19660
rect 32600 19378 32628 19654
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32220 12436 32272 12442
rect 32220 12378 32272 12384
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32128 11756 32180 11762
rect 32128 11698 32180 11704
rect 32140 11082 32168 11698
rect 32232 11558 32260 12378
rect 32312 12232 32364 12238
rect 32312 12174 32364 12180
rect 32324 11694 32352 12174
rect 32312 11688 32364 11694
rect 32312 11630 32364 11636
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 32140 10674 32168 11018
rect 32128 10668 32180 10674
rect 32128 10610 32180 10616
rect 32232 10470 32260 11494
rect 32324 11354 32352 11630
rect 32312 11348 32364 11354
rect 32312 11290 32364 11296
rect 32220 10464 32272 10470
rect 32220 10406 32272 10412
rect 31944 10124 31996 10130
rect 31944 10066 31996 10072
rect 31864 9982 31984 10010
rect 31760 9512 31812 9518
rect 31758 9480 31760 9489
rect 31812 9480 31814 9489
rect 31758 9415 31814 9424
rect 31772 9389 31800 9415
rect 31956 8945 31984 9982
rect 32036 9988 32088 9994
rect 32036 9930 32088 9936
rect 32312 9988 32364 9994
rect 32312 9930 32364 9936
rect 32048 9722 32076 9930
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 32324 9178 32352 9930
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 32416 9353 32444 9590
rect 32402 9344 32458 9353
rect 32402 9279 32458 9288
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32402 9072 32458 9081
rect 32402 9007 32404 9016
rect 32456 9007 32458 9016
rect 32404 8978 32456 8984
rect 31942 8936 31998 8945
rect 31942 8871 31998 8880
rect 32496 8900 32548 8906
rect 32496 8842 32548 8848
rect 32036 8832 32088 8838
rect 32036 8774 32088 8780
rect 32048 8401 32076 8774
rect 32034 8392 32090 8401
rect 32034 8327 32090 8336
rect 31680 4508 31800 4536
rect 31576 4480 31628 4486
rect 31576 4422 31628 4428
rect 31588 3534 31616 4422
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 31576 3392 31628 3398
rect 31576 3334 31628 3340
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 31312 3182 31524 3210
rect 31116 3052 31168 3058
rect 31116 2994 31168 3000
rect 31312 2774 31340 3182
rect 31392 3120 31444 3126
rect 31588 3108 31616 3334
rect 31444 3080 31616 3108
rect 31772 3074 31800 4508
rect 31944 4140 31996 4146
rect 31944 4082 31996 4088
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31864 3097 31892 3130
rect 31392 3062 31444 3068
rect 31680 3046 31800 3074
rect 31850 3088 31906 3097
rect 31312 2746 31524 2774
rect 31496 2514 31524 2746
rect 31484 2508 31536 2514
rect 31484 2450 31536 2456
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 27988 2304 28040 2310
rect 27988 2246 28040 2252
rect 28000 800 28028 2246
rect 28920 800 28948 2382
rect 29460 2304 29512 2310
rect 29460 2246 29512 2252
rect 29472 800 29500 2246
rect 30392 800 30420 2382
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30852 800 30880 2246
rect 31680 2038 31708 3046
rect 31850 3023 31906 3032
rect 31956 2990 31984 4082
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31852 2440 31904 2446
rect 31852 2382 31904 2388
rect 31668 2032 31720 2038
rect 31668 1974 31720 1980
rect 31864 800 31892 2382
rect 32048 2106 32076 8327
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32140 6730 32168 7142
rect 32324 7002 32352 7346
rect 32416 7206 32444 7346
rect 32508 7342 32536 8842
rect 32496 7336 32548 7342
rect 32496 7278 32548 7284
rect 32404 7200 32456 7206
rect 32404 7142 32456 7148
rect 32312 6996 32364 7002
rect 32312 6938 32364 6944
rect 32128 6724 32180 6730
rect 32128 6666 32180 6672
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 32220 6384 32272 6390
rect 32220 6326 32272 6332
rect 32232 5778 32260 6326
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32140 3942 32168 4082
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 32140 3534 32168 3878
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32324 2990 32352 3334
rect 32416 3058 32444 6598
rect 32496 5568 32548 5574
rect 32496 5510 32548 5516
rect 32508 3942 32536 5510
rect 32600 3942 32628 18566
rect 32680 17332 32732 17338
rect 32680 17274 32732 17280
rect 32692 12434 32720 17274
rect 32784 17202 32812 18702
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 32864 16720 32916 16726
rect 32864 16662 32916 16668
rect 32772 15632 32824 15638
rect 32772 15574 32824 15580
rect 32784 14346 32812 15574
rect 32772 14340 32824 14346
rect 32772 14282 32824 14288
rect 32784 14074 32812 14282
rect 32772 14068 32824 14074
rect 32772 14010 32824 14016
rect 32876 13530 32904 16662
rect 33140 16244 33192 16250
rect 33140 16186 33192 16192
rect 33152 16153 33180 16186
rect 33138 16144 33194 16153
rect 33138 16079 33194 16088
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33336 14822 33364 15982
rect 33324 14816 33376 14822
rect 33324 14758 33376 14764
rect 33428 13530 33456 21286
rect 33612 20942 33640 21966
rect 33690 21584 33746 21593
rect 33690 21519 33692 21528
rect 33744 21519 33746 21528
rect 33692 21490 33744 21496
rect 33600 20936 33652 20942
rect 33600 20878 33652 20884
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33520 18329 33548 18770
rect 33506 18320 33562 18329
rect 33506 18255 33508 18264
rect 33560 18255 33562 18264
rect 33508 18226 33560 18232
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33520 15502 33548 15846
rect 33508 15496 33560 15502
rect 33508 15438 33560 15444
rect 33612 14414 33640 20878
rect 34256 20874 34284 22066
rect 34808 22030 34836 22374
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 36280 22098 36308 22374
rect 36268 22092 36320 22098
rect 36268 22034 36320 22040
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34428 21956 34480 21962
rect 34428 21898 34480 21904
rect 34440 21350 34468 21898
rect 35716 21888 35768 21894
rect 35716 21830 35768 21836
rect 35728 21690 35756 21830
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35256 21616 35308 21622
rect 35808 21616 35860 21622
rect 35308 21576 35388 21604
rect 35256 21558 35308 21564
rect 34704 21548 34756 21554
rect 34704 21490 34756 21496
rect 34428 21344 34480 21350
rect 34428 21286 34480 21292
rect 34612 21344 34664 21350
rect 34612 21286 34664 21292
rect 34244 20868 34296 20874
rect 34244 20810 34296 20816
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34072 19514 34100 20538
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 33876 19372 33928 19378
rect 33876 19314 33928 19320
rect 33888 18766 33916 19314
rect 33876 18760 33928 18766
rect 33876 18702 33928 18708
rect 33888 18222 33916 18702
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33968 18148 34020 18154
rect 33968 18090 34020 18096
rect 33692 17604 33744 17610
rect 33692 17546 33744 17552
rect 33704 14906 33732 17546
rect 33980 16590 34008 18090
rect 34060 17604 34112 17610
rect 34060 17546 34112 17552
rect 33784 16584 33836 16590
rect 33784 16526 33836 16532
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 33796 15706 33824 16526
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 33888 16114 33916 16390
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33968 16040 34020 16046
rect 33968 15982 34020 15988
rect 33980 15706 34008 15982
rect 33784 15700 33836 15706
rect 33784 15642 33836 15648
rect 33968 15700 34020 15706
rect 33968 15642 34020 15648
rect 34072 15570 34100 17546
rect 34060 15564 34112 15570
rect 34060 15506 34112 15512
rect 33704 14878 33916 14906
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33888 14278 33916 14878
rect 34072 14618 34100 15506
rect 34060 14612 34112 14618
rect 34060 14554 34112 14560
rect 34060 14476 34112 14482
rect 34060 14418 34112 14424
rect 33876 14272 33928 14278
rect 33876 14214 33928 14220
rect 33690 13968 33746 13977
rect 33690 13903 33692 13912
rect 33744 13903 33746 13912
rect 33692 13874 33744 13880
rect 32864 13524 32916 13530
rect 32864 13466 32916 13472
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 32692 12406 32812 12434
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32692 9586 32720 9862
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32496 3936 32548 3942
rect 32496 3878 32548 3884
rect 32588 3936 32640 3942
rect 32588 3878 32640 3884
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 32036 2100 32088 2106
rect 32036 2042 32088 2048
rect 32324 800 32352 2790
rect 32784 2774 32812 12406
rect 32876 8537 32904 13466
rect 33140 13252 33192 13258
rect 33140 13194 33192 13200
rect 33152 12986 33180 13194
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 32956 11552 33008 11558
rect 32956 11494 33008 11500
rect 33324 11552 33376 11558
rect 33324 11494 33376 11500
rect 32968 11150 32996 11494
rect 33336 11150 33364 11494
rect 32956 11144 33008 11150
rect 32956 11086 33008 11092
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 33048 11008 33100 11014
rect 33048 10950 33100 10956
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33060 10810 33088 10950
rect 33048 10804 33100 10810
rect 33048 10746 33100 10752
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 33152 9586 33180 9930
rect 33244 9674 33272 10950
rect 33336 10418 33364 11086
rect 33428 10538 33456 13466
rect 33704 12102 33732 13874
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33888 11558 33916 14214
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 33980 11830 34008 12174
rect 33968 11824 34020 11830
rect 33968 11766 34020 11772
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33600 11348 33652 11354
rect 33600 11290 33652 11296
rect 33416 10532 33468 10538
rect 33416 10474 33468 10480
rect 33336 10390 33456 10418
rect 33244 9646 33364 9674
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33048 9444 33100 9450
rect 33048 9386 33100 9392
rect 32862 8528 32918 8537
rect 32862 8463 32918 8472
rect 32876 7478 32904 8463
rect 33060 8090 33088 9386
rect 33048 8084 33100 8090
rect 33048 8026 33100 8032
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 33152 7410 33180 9522
rect 33232 7812 33284 7818
rect 33232 7754 33284 7760
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33152 6730 33180 7346
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33060 5302 33088 5782
rect 33152 5642 33180 6666
rect 33244 6662 33272 7754
rect 33336 7206 33364 9646
rect 33428 8294 33456 10390
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33520 9586 33548 9998
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33520 9178 33548 9522
rect 33508 9172 33560 9178
rect 33508 9114 33560 9120
rect 33612 8906 33640 11290
rect 33692 9580 33744 9586
rect 34072 9568 34100 14418
rect 33692 9522 33744 9528
rect 33888 9540 34100 9568
rect 33704 9450 33732 9522
rect 33784 9512 33836 9518
rect 33782 9480 33784 9489
rect 33836 9480 33838 9489
rect 33692 9444 33744 9450
rect 33782 9415 33838 9424
rect 33692 9386 33744 9392
rect 33692 9036 33744 9042
rect 33692 8978 33744 8984
rect 33600 8900 33652 8906
rect 33520 8860 33600 8888
rect 33416 8288 33468 8294
rect 33416 8230 33468 8236
rect 33520 8090 33548 8860
rect 33600 8842 33652 8848
rect 33704 8786 33732 8978
rect 33612 8758 33732 8786
rect 33782 8800 33838 8809
rect 33508 8084 33560 8090
rect 33508 8026 33560 8032
rect 33612 7954 33640 8758
rect 33782 8735 33838 8744
rect 33796 8498 33824 8735
rect 33784 8492 33836 8498
rect 33784 8434 33836 8440
rect 33600 7948 33652 7954
rect 33600 7890 33652 7896
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6458 33364 6598
rect 33324 6452 33376 6458
rect 33324 6394 33376 6400
rect 33416 6316 33468 6322
rect 33416 6258 33468 6264
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 33048 5296 33100 5302
rect 33048 5238 33100 5244
rect 33048 5160 33100 5166
rect 33048 5102 33100 5108
rect 33060 4282 33088 5102
rect 33232 4752 33284 4758
rect 33232 4694 33284 4700
rect 33140 4548 33192 4554
rect 33244 4536 33272 4694
rect 33324 4616 33376 4622
rect 33192 4508 33272 4536
rect 33322 4584 33324 4593
rect 33376 4584 33378 4593
rect 33322 4519 33378 4528
rect 33140 4490 33192 4496
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 33060 4078 33088 4218
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 33428 3058 33456 6258
rect 33692 6180 33744 6186
rect 33692 6122 33744 6128
rect 33598 5264 33654 5273
rect 33598 5199 33654 5208
rect 33508 5024 33560 5030
rect 33508 4966 33560 4972
rect 33520 4622 33548 4966
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 33612 4554 33640 5199
rect 33704 4622 33732 6122
rect 33888 4758 33916 9540
rect 34164 9466 34192 19382
rect 34256 14482 34284 20810
rect 34428 16176 34480 16182
rect 34426 16144 34428 16153
rect 34520 16176 34572 16182
rect 34480 16144 34482 16153
rect 34520 16118 34572 16124
rect 34426 16079 34482 16088
rect 34532 15094 34560 16118
rect 34520 15088 34572 15094
rect 34520 15030 34572 15036
rect 34244 14476 34296 14482
rect 34244 14418 34296 14424
rect 34244 13932 34296 13938
rect 34244 13874 34296 13880
rect 34256 13734 34284 13874
rect 34532 13870 34560 15030
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 34244 13728 34296 13734
rect 34244 13670 34296 13676
rect 34256 13462 34284 13670
rect 34244 13456 34296 13462
rect 34244 13398 34296 13404
rect 34532 12442 34560 13806
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34532 11762 34560 12378
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 34072 9438 34192 9466
rect 33968 8832 34020 8838
rect 33968 8774 34020 8780
rect 33980 8566 34008 8774
rect 33968 8560 34020 8566
rect 33968 8502 34020 8508
rect 33876 4752 33928 4758
rect 33876 4694 33928 4700
rect 33692 4616 33744 4622
rect 33692 4558 33744 4564
rect 33600 4548 33652 4554
rect 33600 4490 33652 4496
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 33784 4140 33836 4146
rect 33784 4082 33836 4088
rect 33796 4010 33824 4082
rect 33784 4004 33836 4010
rect 33784 3946 33836 3952
rect 33876 3120 33928 3126
rect 33980 3108 34008 4422
rect 33928 3080 34008 3108
rect 33876 3062 33928 3068
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 34072 2774 34100 9438
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 34164 8974 34192 9318
rect 34336 9104 34388 9110
rect 34334 9072 34336 9081
rect 34388 9072 34390 9081
rect 34334 9007 34390 9016
rect 34152 8968 34204 8974
rect 34152 8910 34204 8916
rect 34336 8900 34388 8906
rect 34336 8842 34388 8848
rect 34348 8809 34376 8842
rect 34334 8800 34390 8809
rect 34334 8735 34390 8744
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34348 8378 34376 8570
rect 34164 8350 34376 8378
rect 34164 8294 34192 8350
rect 34152 8288 34204 8294
rect 34152 8230 34204 8236
rect 34244 8288 34296 8294
rect 34296 8236 34376 8242
rect 34244 8230 34376 8236
rect 34256 8214 34376 8230
rect 34348 7750 34376 8214
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 34152 6724 34204 6730
rect 34152 6666 34204 6672
rect 34164 6322 34192 6666
rect 34152 6316 34204 6322
rect 34152 6258 34204 6264
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 5030 34284 6258
rect 34348 5234 34376 7686
rect 34428 6112 34480 6118
rect 34428 6054 34480 6060
rect 34440 5370 34468 6054
rect 34428 5364 34480 5370
rect 34428 5306 34480 5312
rect 34336 5228 34388 5234
rect 34336 5170 34388 5176
rect 34244 5024 34296 5030
rect 34244 4966 34296 4972
rect 34244 4684 34296 4690
rect 34244 4626 34296 4632
rect 34256 4486 34284 4626
rect 34244 4480 34296 4486
rect 34244 4422 34296 4428
rect 32784 2746 32996 2774
rect 32968 2582 32996 2746
rect 33520 2746 34100 2774
rect 34348 2774 34376 5170
rect 34440 3466 34468 5306
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34532 3058 34560 3334
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 34348 2746 34468 2774
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 33336 800 33364 2450
rect 33520 1494 33548 2746
rect 34440 2446 34468 2746
rect 34624 2650 34652 21286
rect 34716 20942 34744 21490
rect 34796 21412 34848 21418
rect 34796 21354 34848 21360
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34808 20806 34836 21354
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 20874 35388 21576
rect 35806 21584 35808 21593
rect 35860 21584 35862 21593
rect 35440 21548 35492 21554
rect 35806 21519 35862 21528
rect 36176 21548 36228 21554
rect 35440 21490 35492 21496
rect 36176 21490 36228 21496
rect 35452 21350 35480 21490
rect 35532 21412 35584 21418
rect 35532 21354 35584 21360
rect 35808 21412 35860 21418
rect 35808 21354 35860 21360
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35348 20868 35400 20874
rect 35348 20810 35400 20816
rect 35440 20868 35492 20874
rect 35440 20810 35492 20816
rect 34796 20800 34848 20806
rect 34796 20742 34848 20748
rect 35360 20534 35388 20810
rect 35348 20528 35400 20534
rect 35348 20470 35400 20476
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34808 19786 34836 20402
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34796 19780 34848 19786
rect 34796 19722 34848 19728
rect 34808 19310 34836 19722
rect 35360 19378 35388 20470
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34808 17678 34836 18158
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34716 12170 34744 17478
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34808 15502 34836 16458
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34808 13530 34836 13874
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 34796 13388 34848 13394
rect 34796 13330 34848 13336
rect 34704 12164 34756 12170
rect 34704 12106 34756 12112
rect 34808 10266 34836 13330
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35360 11354 35388 11698
rect 35348 11348 35400 11354
rect 35348 11290 35400 11296
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34704 10056 34756 10062
rect 34704 9998 34756 10004
rect 34716 8838 34744 9998
rect 35256 9920 35308 9926
rect 35256 9862 35308 9868
rect 35268 9450 35296 9862
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 35348 9376 35400 9382
rect 35348 9318 35400 9324
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 35360 8974 35388 9318
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 34704 8832 34756 8838
rect 34704 8774 34756 8780
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35452 7562 35480 20810
rect 35544 16454 35572 21354
rect 35820 21078 35848 21354
rect 35808 21072 35860 21078
rect 35808 21014 35860 21020
rect 35808 20936 35860 20942
rect 35808 20878 35860 20884
rect 35820 20806 35848 20878
rect 36188 20806 36216 21490
rect 36280 20942 36308 22034
rect 39120 22024 39172 22030
rect 39120 21966 39172 21972
rect 37832 21956 37884 21962
rect 37832 21898 37884 21904
rect 38292 21956 38344 21962
rect 38292 21898 38344 21904
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 37844 20874 37872 21898
rect 38016 21412 38068 21418
rect 38016 21354 38068 21360
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 36544 20868 36596 20874
rect 36544 20810 36596 20816
rect 37832 20868 37884 20874
rect 37832 20810 37884 20816
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 35716 20460 35768 20466
rect 35820 20448 35848 20742
rect 36188 20466 36216 20742
rect 36372 20602 36400 20810
rect 36360 20596 36412 20602
rect 36360 20538 36412 20544
rect 36452 20528 36504 20534
rect 36452 20470 36504 20476
rect 35768 20420 35848 20448
rect 35716 20402 35768 20408
rect 35820 19854 35848 20420
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 35808 19848 35860 19854
rect 35808 19790 35860 19796
rect 36188 19802 36216 20402
rect 36268 19848 36320 19854
rect 36188 19796 36268 19802
rect 36188 19790 36320 19796
rect 35820 18290 35848 19790
rect 36084 19780 36136 19786
rect 36084 19722 36136 19728
rect 36188 19774 36308 19790
rect 36096 19174 36124 19722
rect 36084 19168 36136 19174
rect 36084 19110 36136 19116
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 36004 18290 36032 18702
rect 36096 18630 36124 19110
rect 36188 18902 36216 19774
rect 36176 18896 36228 18902
rect 36176 18838 36228 18844
rect 36084 18624 36136 18630
rect 36084 18566 36136 18572
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 36004 17542 36032 18226
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 35624 16788 35676 16794
rect 35624 16730 35676 16736
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35532 11552 35584 11558
rect 35532 11494 35584 11500
rect 35544 11354 35572 11494
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35532 10736 35584 10742
rect 35532 10678 35584 10684
rect 35544 9586 35572 10678
rect 35636 9926 35664 16730
rect 35992 16516 36044 16522
rect 35992 16458 36044 16464
rect 36004 15502 36032 16458
rect 36268 15632 36320 15638
rect 36268 15574 36320 15580
rect 35992 15496 36044 15502
rect 35992 15438 36044 15444
rect 36004 15026 36032 15438
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 35900 14612 35952 14618
rect 35900 14554 35952 14560
rect 35808 14340 35860 14346
rect 35808 14282 35860 14288
rect 35716 11348 35768 11354
rect 35716 11290 35768 11296
rect 35728 11150 35756 11290
rect 35716 11144 35768 11150
rect 35716 11086 35768 11092
rect 35624 9920 35676 9926
rect 35624 9862 35676 9868
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35532 9444 35584 9450
rect 35532 9386 35584 9392
rect 35544 9217 35572 9386
rect 35530 9208 35586 9217
rect 35530 9143 35586 9152
rect 35452 7534 35664 7562
rect 35440 7404 35492 7410
rect 35440 7346 35492 7352
rect 35348 7268 35400 7274
rect 35348 7210 35400 7216
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35360 6662 35388 7210
rect 35452 6730 35480 7346
rect 35440 6724 35492 6730
rect 35440 6666 35492 6672
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 35360 6322 35388 6598
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34704 6112 34756 6118
rect 34704 6054 34756 6060
rect 34716 5846 34744 6054
rect 34704 5840 34756 5846
rect 34702 5808 34704 5817
rect 34808 5828 34836 6190
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35532 5840 35584 5846
rect 34756 5808 34758 5817
rect 34808 5800 35204 5828
rect 34702 5743 34758 5752
rect 34704 5704 34756 5710
rect 34704 5646 34756 5652
rect 34716 3194 34744 5646
rect 35176 5642 35204 5800
rect 35532 5782 35584 5788
rect 35164 5636 35216 5642
rect 35164 5578 35216 5584
rect 35440 5568 35492 5574
rect 35440 5510 35492 5516
rect 35348 5296 35400 5302
rect 35452 5284 35480 5510
rect 35400 5256 35480 5284
rect 35348 5238 35400 5244
rect 35256 5092 35308 5098
rect 35308 5052 35388 5080
rect 35256 5034 35308 5040
rect 35360 5001 35388 5052
rect 35346 4992 35402 5001
rect 34934 4924 35242 4944
rect 35346 4927 35402 4936
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35254 4720 35310 4729
rect 35254 4655 35310 4664
rect 35268 4622 35296 4655
rect 35452 4622 35480 5256
rect 35544 4826 35572 5782
rect 35532 4820 35584 4826
rect 35532 4762 35584 4768
rect 35256 4616 35308 4622
rect 35256 4558 35308 4564
rect 35440 4616 35492 4622
rect 35440 4558 35492 4564
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35360 3534 35388 3878
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 34716 2378 34744 3130
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 33784 2304 33836 2310
rect 33784 2246 33836 2252
rect 33508 1488 33560 1494
rect 33508 1430 33560 1436
rect 33796 800 33824 2246
rect 34808 800 34836 3470
rect 35544 3466 35572 4762
rect 35532 3460 35584 3466
rect 35532 3402 35584 3408
rect 35256 2984 35308 2990
rect 35254 2952 35256 2961
rect 35308 2952 35310 2961
rect 35254 2887 35310 2896
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35636 2650 35664 7534
rect 35728 4729 35756 11086
rect 35820 8566 35848 14282
rect 35912 13938 35940 14554
rect 35900 13932 35952 13938
rect 35900 13874 35952 13880
rect 35912 13734 35940 13874
rect 35900 13728 35952 13734
rect 35900 13670 35952 13676
rect 35912 13258 35940 13670
rect 35900 13252 35952 13258
rect 35900 13194 35952 13200
rect 36004 11830 36032 14962
rect 36176 14272 36228 14278
rect 36176 14214 36228 14220
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 36096 12442 36124 13262
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 35992 11824 36044 11830
rect 35992 11766 36044 11772
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 35912 9489 35940 10406
rect 35898 9480 35954 9489
rect 35898 9415 35954 9424
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35808 8424 35860 8430
rect 35806 8392 35808 8401
rect 35860 8392 35862 8401
rect 35806 8327 35862 8336
rect 35806 5808 35862 5817
rect 35806 5743 35862 5752
rect 35714 4720 35770 4729
rect 35714 4655 35770 4664
rect 35716 4616 35768 4622
rect 35820 4604 35848 5743
rect 35912 5642 35940 8978
rect 36004 7206 36032 11766
rect 36096 11558 36124 12378
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 36084 11008 36136 11014
rect 36084 10950 36136 10956
rect 36096 10674 36124 10950
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 35992 7200 36044 7206
rect 35992 7142 36044 7148
rect 36004 7002 36032 7142
rect 35992 6996 36044 7002
rect 35992 6938 36044 6944
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 36004 6254 36032 6666
rect 36096 6458 36124 10202
rect 36188 9994 36216 14214
rect 36280 13326 36308 15574
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 36372 13530 36400 14350
rect 36360 13524 36412 13530
rect 36360 13466 36412 13472
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 36360 11620 36412 11626
rect 36360 11562 36412 11568
rect 36372 11150 36400 11562
rect 36268 11144 36320 11150
rect 36268 11086 36320 11092
rect 36360 11144 36412 11150
rect 36360 11086 36412 11092
rect 36280 10996 36308 11086
rect 36360 11008 36412 11014
rect 36280 10968 36360 10996
rect 36360 10950 36412 10956
rect 36372 10674 36400 10950
rect 36360 10668 36412 10674
rect 36360 10610 36412 10616
rect 36176 9988 36228 9994
rect 36176 9930 36228 9936
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 36280 9586 36308 9862
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36176 9376 36228 9382
rect 36176 9318 36228 9324
rect 36188 8498 36216 9318
rect 36280 8498 36308 9522
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 36360 8288 36412 8294
rect 36360 8230 36412 8236
rect 36188 7886 36216 8230
rect 36372 7886 36400 8230
rect 36176 7880 36228 7886
rect 36360 7880 36412 7886
rect 36228 7840 36308 7868
rect 36176 7822 36228 7828
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 36188 7002 36216 7142
rect 36176 6996 36228 7002
rect 36176 6938 36228 6944
rect 36280 6458 36308 7840
rect 36360 7822 36412 7828
rect 36372 7546 36400 7822
rect 36360 7540 36412 7546
rect 36360 7482 36412 7488
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 36372 6322 36400 7482
rect 36464 7478 36492 20470
rect 36556 16674 36584 20810
rect 38028 19854 38056 21354
rect 38304 21146 38332 21898
rect 38660 21888 38712 21894
rect 38660 21830 38712 21836
rect 38672 21554 38700 21830
rect 38660 21548 38712 21554
rect 38660 21490 38712 21496
rect 38292 21140 38344 21146
rect 38292 21082 38344 21088
rect 38200 20392 38252 20398
rect 38200 20334 38252 20340
rect 38016 19848 38068 19854
rect 38016 19790 38068 19796
rect 37096 19780 37148 19786
rect 37096 19722 37148 19728
rect 37004 19168 37056 19174
rect 37004 19110 37056 19116
rect 36636 18964 36688 18970
rect 36636 18906 36688 18912
rect 36648 18766 36676 18906
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 37016 18698 37044 19110
rect 36912 18692 36964 18698
rect 36912 18634 36964 18640
rect 37004 18692 37056 18698
rect 37004 18634 37056 18640
rect 36636 18624 36688 18630
rect 36636 18566 36688 18572
rect 36648 18465 36676 18566
rect 36634 18456 36690 18465
rect 36634 18391 36690 18400
rect 36556 16646 36676 16674
rect 36544 13796 36596 13802
rect 36544 13738 36596 13744
rect 36556 12238 36584 13738
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36544 11144 36596 11150
rect 36544 11086 36596 11092
rect 36556 10130 36584 11086
rect 36544 10124 36596 10130
rect 36544 10066 36596 10072
rect 36544 8832 36596 8838
rect 36544 8774 36596 8780
rect 36556 8634 36584 8774
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36648 7562 36676 16646
rect 36728 15156 36780 15162
rect 36728 15098 36780 15104
rect 36740 14414 36768 15098
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 36740 13938 36768 14350
rect 36728 13932 36780 13938
rect 36728 13874 36780 13880
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36740 10266 36768 13466
rect 36820 13456 36872 13462
rect 36820 13398 36872 13404
rect 36924 13410 36952 18634
rect 37004 16652 37056 16658
rect 37004 16594 37056 16600
rect 37016 14958 37044 16594
rect 37004 14952 37056 14958
rect 37004 14894 37056 14900
rect 37004 14408 37056 14414
rect 37004 14350 37056 14356
rect 37016 13530 37044 14350
rect 37004 13524 37056 13530
rect 37004 13466 37056 13472
rect 36728 10260 36780 10266
rect 36728 10202 36780 10208
rect 36832 9489 36860 13398
rect 36924 13382 37044 13410
rect 36912 13320 36964 13326
rect 36912 13262 36964 13268
rect 36818 9480 36874 9489
rect 36818 9415 36874 9424
rect 36832 9042 36860 9415
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36544 7540 36596 7546
rect 36648 7534 36860 7562
rect 36544 7482 36596 7488
rect 36452 7472 36504 7478
rect 36452 7414 36504 7420
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 36372 5710 36400 6258
rect 36360 5704 36412 5710
rect 36360 5646 36412 5652
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35992 5364 36044 5370
rect 35992 5306 36044 5312
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35900 5024 35952 5030
rect 35900 4966 35952 4972
rect 35912 4622 35940 4966
rect 36004 4826 36032 5306
rect 36096 5273 36124 5306
rect 36082 5264 36138 5273
rect 36082 5199 36138 5208
rect 36082 4992 36138 5001
rect 36082 4927 36138 4936
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 36096 4690 36124 4927
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 35768 4576 35848 4604
rect 35716 4558 35768 4564
rect 35820 4010 35848 4576
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35912 4078 35940 4558
rect 36084 4208 36136 4214
rect 36084 4150 36136 4156
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 35808 4004 35860 4010
rect 35808 3946 35860 3952
rect 35912 3738 35940 4014
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 36096 3534 36124 4150
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36464 3602 36492 3878
rect 36446 3596 36498 3602
rect 36446 3538 36498 3544
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 35624 2644 35676 2650
rect 35624 2586 35676 2592
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 35256 2304 35308 2310
rect 35256 2246 35308 2252
rect 35268 800 35296 2246
rect 36280 800 36308 2382
rect 36556 2310 36584 7482
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 36740 5642 36768 6054
rect 36728 5636 36780 5642
rect 36728 5578 36780 5584
rect 36636 4004 36688 4010
rect 36636 3946 36688 3952
rect 36648 3534 36676 3946
rect 36728 3664 36780 3670
rect 36728 3606 36780 3612
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 36740 3233 36768 3606
rect 36726 3224 36782 3233
rect 36726 3159 36782 3168
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 36544 2304 36596 2310
rect 36544 2246 36596 2252
rect 36740 800 36768 2790
rect 36832 2774 36860 7534
rect 36924 6322 36952 13262
rect 37016 7546 37044 13382
rect 37108 12434 37136 19722
rect 38028 19242 38056 19790
rect 38212 19786 38240 20334
rect 38292 19848 38344 19854
rect 38292 19790 38344 19796
rect 38200 19780 38252 19786
rect 38200 19722 38252 19728
rect 38212 19310 38240 19722
rect 38304 19378 38332 19790
rect 38292 19372 38344 19378
rect 38292 19314 38344 19320
rect 38200 19304 38252 19310
rect 38200 19246 38252 19252
rect 38016 19236 38068 19242
rect 38016 19178 38068 19184
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37372 18760 37424 18766
rect 37372 18702 37424 18708
rect 37200 18290 37228 18702
rect 37384 18358 37412 18702
rect 37556 18692 37608 18698
rect 37556 18634 37608 18640
rect 37372 18352 37424 18358
rect 37372 18294 37424 18300
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37372 18080 37424 18086
rect 37372 18022 37424 18028
rect 37384 17678 37412 18022
rect 37476 17882 37504 18226
rect 37464 17876 37516 17882
rect 37464 17818 37516 17824
rect 37372 17672 37424 17678
rect 37372 17614 37424 17620
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 37200 16658 37228 17478
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 37292 16454 37320 17138
rect 37372 17128 37424 17134
rect 37372 17070 37424 17076
rect 37384 16658 37412 17070
rect 37372 16652 37424 16658
rect 37372 16594 37424 16600
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 37384 16266 37412 16594
rect 37292 16238 37412 16266
rect 37292 15094 37320 16238
rect 37372 15632 37424 15638
rect 37372 15574 37424 15580
rect 37280 15088 37332 15094
rect 37280 15030 37332 15036
rect 37384 14618 37412 15574
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37476 14618 37504 14962
rect 37372 14612 37424 14618
rect 37372 14554 37424 14560
rect 37464 14612 37516 14618
rect 37464 14554 37516 14560
rect 37280 12640 37332 12646
rect 37280 12582 37332 12588
rect 37108 12406 37228 12434
rect 37096 12232 37148 12238
rect 37096 12174 37148 12180
rect 37108 11762 37136 12174
rect 37096 11756 37148 11762
rect 37096 11698 37148 11704
rect 37004 7540 37056 7546
rect 37004 7482 37056 7488
rect 37096 7472 37148 7478
rect 37096 7414 37148 7420
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 37016 6934 37044 7210
rect 37004 6928 37056 6934
rect 37004 6870 37056 6876
rect 37016 6798 37044 6870
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 36912 6316 36964 6322
rect 36912 6258 36964 6264
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 36924 3126 36952 3674
rect 37004 3528 37056 3534
rect 37004 3470 37056 3476
rect 36912 3120 36964 3126
rect 36912 3062 36964 3068
rect 37016 2922 37044 3470
rect 37004 2916 37056 2922
rect 37004 2858 37056 2864
rect 36832 2746 37044 2774
rect 37016 2582 37044 2746
rect 37004 2576 37056 2582
rect 37004 2518 37056 2524
rect 37108 2378 37136 7414
rect 37096 2372 37148 2378
rect 37096 2314 37148 2320
rect 37200 2106 37228 12406
rect 37292 12238 37320 12582
rect 37568 12434 37596 18634
rect 38028 18630 38056 19178
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 37844 18426 37872 18566
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 38028 18222 38056 18566
rect 38212 18222 38240 19246
rect 38672 18902 38700 21490
rect 38844 21480 38896 21486
rect 38844 21422 38896 21428
rect 38752 21344 38804 21350
rect 38752 21286 38804 21292
rect 38764 20942 38792 21286
rect 38752 20936 38804 20942
rect 38752 20878 38804 20884
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38764 20058 38792 20402
rect 38752 20052 38804 20058
rect 38752 19994 38804 20000
rect 38856 19922 38884 21422
rect 39132 20398 39160 21966
rect 39856 20868 39908 20874
rect 39856 20810 39908 20816
rect 39120 20392 39172 20398
rect 39120 20334 39172 20340
rect 39132 20058 39160 20334
rect 39120 20052 39172 20058
rect 39120 19994 39172 20000
rect 38844 19916 38896 19922
rect 38844 19858 38896 19864
rect 39120 19916 39172 19922
rect 39120 19858 39172 19864
rect 39028 19848 39080 19854
rect 39028 19790 39080 19796
rect 39040 19514 39068 19790
rect 39132 19718 39160 19858
rect 39120 19712 39172 19718
rect 39120 19654 39172 19660
rect 39028 19508 39080 19514
rect 39028 19450 39080 19456
rect 38660 18896 38712 18902
rect 38660 18838 38712 18844
rect 38936 18352 38988 18358
rect 38936 18294 38988 18300
rect 38016 18216 38068 18222
rect 38016 18158 38068 18164
rect 38200 18216 38252 18222
rect 38200 18158 38252 18164
rect 38028 17746 38056 18158
rect 38016 17740 38068 17746
rect 38016 17682 38068 17688
rect 38948 17338 38976 18294
rect 38936 17332 38988 17338
rect 38936 17274 38988 17280
rect 38660 15564 38712 15570
rect 38660 15506 38712 15512
rect 37924 15496 37976 15502
rect 37924 15438 37976 15444
rect 37648 15428 37700 15434
rect 37648 15370 37700 15376
rect 37660 15162 37688 15370
rect 37832 15360 37884 15366
rect 37832 15302 37884 15308
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37844 14278 37872 15302
rect 37936 14482 37964 15438
rect 38672 14618 38700 15506
rect 38752 15020 38804 15026
rect 38752 14962 38804 14968
rect 38660 14612 38712 14618
rect 38660 14554 38712 14560
rect 37924 14476 37976 14482
rect 37924 14418 37976 14424
rect 38476 14476 38528 14482
rect 38476 14418 38528 14424
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37568 12406 37688 12434
rect 37280 12232 37332 12238
rect 37280 12174 37332 12180
rect 37292 6798 37320 12174
rect 37372 12096 37424 12102
rect 37372 12038 37424 12044
rect 37464 12096 37516 12102
rect 37464 12038 37516 12044
rect 37384 11830 37412 12038
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 37476 10062 37504 12038
rect 37556 11552 37608 11558
rect 37556 11494 37608 11500
rect 37568 11218 37596 11494
rect 37556 11212 37608 11218
rect 37556 11154 37608 11160
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37476 7478 37504 9998
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 37568 9178 37596 9318
rect 37556 9172 37608 9178
rect 37556 9114 37608 9120
rect 37464 7472 37516 7478
rect 37464 7414 37516 7420
rect 37372 6928 37424 6934
rect 37372 6870 37424 6876
rect 37280 6792 37332 6798
rect 37280 6734 37332 6740
rect 37384 6497 37412 6870
rect 37556 6860 37608 6866
rect 37556 6802 37608 6808
rect 37370 6488 37426 6497
rect 37370 6423 37426 6432
rect 37464 4752 37516 4758
rect 37464 4694 37516 4700
rect 37476 4282 37504 4694
rect 37568 4622 37596 6802
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37568 4486 37596 4558
rect 37556 4480 37608 4486
rect 37556 4422 37608 4428
rect 37464 4276 37516 4282
rect 37464 4218 37516 4224
rect 37556 2440 37608 2446
rect 37556 2382 37608 2388
rect 37188 2100 37240 2106
rect 37188 2042 37240 2048
rect 37568 2038 37596 2382
rect 37556 2032 37608 2038
rect 37556 1974 37608 1980
rect 37660 1562 37688 12406
rect 38488 12170 38516 14418
rect 38764 13870 38792 14962
rect 39132 14550 39160 19654
rect 39868 17542 39896 20810
rect 40040 20256 40092 20262
rect 40040 20198 40092 20204
rect 40052 19446 40080 20198
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 40040 19440 40092 19446
rect 40040 19382 40092 19388
rect 40052 18766 40080 19382
rect 40040 18760 40092 18766
rect 40040 18702 40092 18708
rect 39948 18692 40000 18698
rect 39948 18634 40000 18640
rect 39960 18358 39988 18634
rect 40408 18624 40460 18630
rect 40408 18566 40460 18572
rect 39948 18352 40000 18358
rect 39948 18294 40000 18300
rect 40040 18284 40092 18290
rect 40040 18226 40092 18232
rect 40052 17882 40080 18226
rect 40420 18222 40448 18566
rect 40512 18222 40540 19994
rect 40408 18216 40460 18222
rect 40408 18158 40460 18164
rect 40500 18216 40552 18222
rect 40500 18158 40552 18164
rect 40316 18080 40368 18086
rect 40316 18022 40368 18028
rect 40040 17876 40092 17882
rect 40040 17818 40092 17824
rect 40328 17678 40356 18022
rect 40512 17746 40540 18158
rect 40500 17740 40552 17746
rect 40500 17682 40552 17688
rect 41052 17740 41104 17746
rect 41052 17682 41104 17688
rect 40040 17672 40092 17678
rect 40040 17614 40092 17620
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 39856 17536 39908 17542
rect 39856 17478 39908 17484
rect 40052 16998 40080 17614
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40052 15722 40080 16934
rect 40224 16652 40276 16658
rect 40224 16594 40276 16600
rect 40236 16114 40264 16594
rect 40592 16584 40644 16590
rect 40592 16526 40644 16532
rect 40316 16516 40368 16522
rect 40316 16458 40368 16464
rect 40224 16108 40276 16114
rect 40224 16050 40276 16056
rect 40052 15694 40172 15722
rect 39120 14544 39172 14550
rect 39120 14486 39172 14492
rect 38752 13864 38804 13870
rect 38752 13806 38804 13812
rect 40040 13864 40092 13870
rect 40040 13806 40092 13812
rect 38764 12850 38792 13806
rect 39764 13320 39816 13326
rect 39764 13262 39816 13268
rect 39776 12850 39804 13262
rect 38752 12844 38804 12850
rect 38752 12786 38804 12792
rect 39764 12844 39816 12850
rect 39764 12786 39816 12792
rect 39212 12708 39264 12714
rect 39212 12650 39264 12656
rect 38476 12164 38528 12170
rect 38476 12106 38528 12112
rect 38384 11688 38436 11694
rect 38384 11630 38436 11636
rect 37740 11552 37792 11558
rect 37740 11494 37792 11500
rect 37752 6390 37780 11494
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 37832 9580 37884 9586
rect 37832 9522 37884 9528
rect 37844 8401 37872 9522
rect 38028 8974 38056 9862
rect 38108 9512 38160 9518
rect 38108 9454 38160 9460
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 37830 8392 37886 8401
rect 37830 8327 37886 8336
rect 37844 7206 37872 8327
rect 37832 7200 37884 7206
rect 37832 7142 37884 7148
rect 37740 6384 37792 6390
rect 37740 6326 37792 6332
rect 37738 4584 37794 4593
rect 37738 4519 37794 4528
rect 37752 4486 37780 4519
rect 37740 4480 37792 4486
rect 37740 4422 37792 4428
rect 37844 4146 37872 7142
rect 37936 5166 37964 8910
rect 38120 8634 38148 9454
rect 38200 9444 38252 9450
rect 38200 9386 38252 9392
rect 38212 8945 38240 9386
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 38396 7886 38424 11630
rect 38488 11150 38516 12106
rect 39224 11762 39252 12650
rect 39856 12640 39908 12646
rect 39856 12582 39908 12588
rect 39868 12238 39896 12582
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 39868 11762 39896 12174
rect 39212 11756 39264 11762
rect 39212 11698 39264 11704
rect 39856 11756 39908 11762
rect 39856 11698 39908 11704
rect 38752 11348 38804 11354
rect 38752 11290 38804 11296
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 38764 10810 38792 11290
rect 38752 10804 38804 10810
rect 38752 10746 38804 10752
rect 39212 10056 39264 10062
rect 39212 9998 39264 10004
rect 39224 9722 39252 9998
rect 38660 9716 38712 9722
rect 38660 9658 38712 9664
rect 39212 9716 39264 9722
rect 39212 9658 39264 9664
rect 38672 8294 38700 9658
rect 38936 9512 38988 9518
rect 38936 9454 38988 9460
rect 39210 9480 39266 9489
rect 38948 9217 38976 9454
rect 39210 9415 39212 9424
rect 39264 9415 39266 9424
rect 39212 9386 39264 9392
rect 38934 9208 38990 9217
rect 40052 9178 40080 13806
rect 38934 9143 38990 9152
rect 40040 9172 40092 9178
rect 40040 9114 40092 9120
rect 39120 9104 39172 9110
rect 39120 9046 39172 9052
rect 39132 8430 39160 9046
rect 39304 8832 39356 8838
rect 39304 8774 39356 8780
rect 39396 8832 39448 8838
rect 39396 8774 39448 8780
rect 39316 8498 39344 8774
rect 39408 8634 39436 8774
rect 40144 8650 40172 15694
rect 40328 14006 40356 16458
rect 40604 15706 40632 16526
rect 40960 16448 41012 16454
rect 40960 16390 41012 16396
rect 40972 16182 41000 16390
rect 40960 16176 41012 16182
rect 40960 16118 41012 16124
rect 41064 16114 41092 17682
rect 42892 17604 42944 17610
rect 42892 17546 42944 17552
rect 42904 17338 42932 17546
rect 42892 17332 42944 17338
rect 42892 17274 42944 17280
rect 43076 17196 43128 17202
rect 43076 17138 43128 17144
rect 43088 16794 43116 17138
rect 43076 16788 43128 16794
rect 43076 16730 43128 16736
rect 43260 16652 43312 16658
rect 43260 16594 43312 16600
rect 41236 16516 41288 16522
rect 41236 16458 41288 16464
rect 41144 16244 41196 16250
rect 41144 16186 41196 16192
rect 41052 16108 41104 16114
rect 41052 16050 41104 16056
rect 40592 15700 40644 15706
rect 40592 15642 40644 15648
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40880 15094 40908 15438
rect 40868 15088 40920 15094
rect 40868 15030 40920 15036
rect 40880 14414 40908 15030
rect 41064 14906 41092 16050
rect 41156 15042 41184 16186
rect 41248 15366 41276 16458
rect 41696 15904 41748 15910
rect 41696 15846 41748 15852
rect 41972 15904 42024 15910
rect 41972 15846 42024 15852
rect 41708 15638 41736 15846
rect 41696 15632 41748 15638
rect 41696 15574 41748 15580
rect 41984 15570 42012 15846
rect 43272 15570 43300 16594
rect 43456 16574 43484 39238
rect 50294 39196 50602 39216
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39120 50602 39140
rect 50294 38108 50602 38128
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38032 50602 38052
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 48320 19712 48372 19718
rect 48320 19654 48372 19660
rect 48332 17882 48360 19654
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 48320 17876 48372 17882
rect 48320 17818 48372 17824
rect 48596 17876 48648 17882
rect 48596 17818 48648 17824
rect 45284 17604 45336 17610
rect 45284 17546 45336 17552
rect 47860 17604 47912 17610
rect 47860 17546 47912 17552
rect 43996 17536 44048 17542
rect 43996 17478 44048 17484
rect 44008 16658 44036 17478
rect 45296 17338 45324 17546
rect 47124 17536 47176 17542
rect 47124 17478 47176 17484
rect 45284 17332 45336 17338
rect 45284 17274 45336 17280
rect 45560 17196 45612 17202
rect 45560 17138 45612 17144
rect 45572 16794 45600 17138
rect 45560 16788 45612 16794
rect 45560 16730 45612 16736
rect 43996 16652 44048 16658
rect 43996 16594 44048 16600
rect 45008 16652 45060 16658
rect 45008 16594 45060 16600
rect 45468 16652 45520 16658
rect 45468 16594 45520 16600
rect 43720 16584 43772 16590
rect 43456 16546 43576 16574
rect 41972 15564 42024 15570
rect 41972 15506 42024 15512
rect 43260 15564 43312 15570
rect 43260 15506 43312 15512
rect 41236 15360 41288 15366
rect 41236 15302 41288 15308
rect 41248 15162 41276 15302
rect 41236 15156 41288 15162
rect 41236 15098 41288 15104
rect 41156 15014 41276 15042
rect 41064 14878 41184 14906
rect 40868 14408 40920 14414
rect 40868 14350 40920 14356
rect 40316 14000 40368 14006
rect 40316 13942 40368 13948
rect 40408 14000 40460 14006
rect 40408 13942 40460 13948
rect 40420 13190 40448 13942
rect 40684 13320 40736 13326
rect 40684 13262 40736 13268
rect 40408 13184 40460 13190
rect 40408 13126 40460 13132
rect 40420 12918 40448 13126
rect 40408 12912 40460 12918
rect 40408 12854 40460 12860
rect 40316 12436 40368 12442
rect 40316 12378 40368 12384
rect 40328 11762 40356 12378
rect 40696 12238 40724 13262
rect 40880 12782 40908 14350
rect 41052 14272 41104 14278
rect 41052 14214 41104 14220
rect 41064 13938 41092 14214
rect 41052 13932 41104 13938
rect 41052 13874 41104 13880
rect 40960 13184 41012 13190
rect 40960 13126 41012 13132
rect 40972 12850 41000 13126
rect 40960 12844 41012 12850
rect 40960 12786 41012 12792
rect 40868 12776 40920 12782
rect 40868 12718 40920 12724
rect 40684 12232 40736 12238
rect 40682 12200 40684 12209
rect 40736 12200 40738 12209
rect 40880 12170 40908 12718
rect 40682 12135 40738 12144
rect 40868 12164 40920 12170
rect 40868 12106 40920 12112
rect 40224 11756 40276 11762
rect 40224 11698 40276 11704
rect 40316 11756 40368 11762
rect 40316 11698 40368 11704
rect 40236 11354 40264 11698
rect 40224 11348 40276 11354
rect 40224 11290 40276 11296
rect 40880 11218 40908 12106
rect 41064 11694 41092 13874
rect 41156 13394 41184 14878
rect 41144 13388 41196 13394
rect 41144 13330 41196 13336
rect 41156 12102 41184 13330
rect 41144 12096 41196 12102
rect 41144 12038 41196 12044
rect 41142 11792 41198 11801
rect 41142 11727 41198 11736
rect 41156 11694 41184 11727
rect 41052 11688 41104 11694
rect 41052 11630 41104 11636
rect 41144 11688 41196 11694
rect 41144 11630 41196 11636
rect 40868 11212 40920 11218
rect 40868 11154 40920 11160
rect 40960 10056 41012 10062
rect 40960 9998 41012 10004
rect 40972 9586 41000 9998
rect 41248 9654 41276 15014
rect 43272 14822 43300 15506
rect 43444 15496 43496 15502
rect 43444 15438 43496 15444
rect 43260 14816 43312 14822
rect 43260 14758 43312 14764
rect 43272 14482 43300 14758
rect 43456 14618 43484 15438
rect 43444 14612 43496 14618
rect 43444 14554 43496 14560
rect 43260 14476 43312 14482
rect 43260 14418 43312 14424
rect 41420 13864 41472 13870
rect 41420 13806 41472 13812
rect 41432 13326 41460 13806
rect 41420 13320 41472 13326
rect 41420 13262 41472 13268
rect 42432 12300 42484 12306
rect 42432 12242 42484 12248
rect 42444 12102 42472 12242
rect 43260 12164 43312 12170
rect 43260 12106 43312 12112
rect 42432 12096 42484 12102
rect 42432 12038 42484 12044
rect 41493 11756 41545 11762
rect 41972 11756 42024 11762
rect 41545 11704 41552 11744
rect 41493 11698 41552 11704
rect 41972 11698 42024 11704
rect 41524 11150 41552 11698
rect 41512 11144 41564 11150
rect 41512 11086 41564 11092
rect 41984 10810 42012 11698
rect 42444 11694 42472 12038
rect 42522 11792 42578 11801
rect 42522 11727 42524 11736
rect 42576 11727 42578 11736
rect 42524 11698 42576 11704
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 42444 11082 42472 11630
rect 43272 11286 43300 12106
rect 43260 11280 43312 11286
rect 43260 11222 43312 11228
rect 42432 11076 42484 11082
rect 42432 11018 42484 11024
rect 42984 11008 43036 11014
rect 42984 10950 43036 10956
rect 41972 10804 42024 10810
rect 41972 10746 42024 10752
rect 42340 10668 42392 10674
rect 42340 10610 42392 10616
rect 42352 10266 42380 10610
rect 42340 10260 42392 10266
rect 42340 10202 42392 10208
rect 42996 10130 43024 10950
rect 43076 10464 43128 10470
rect 43076 10406 43128 10412
rect 42984 10124 43036 10130
rect 42984 10066 43036 10072
rect 43088 10062 43116 10406
rect 41328 10056 41380 10062
rect 41328 9998 41380 10004
rect 41972 10056 42024 10062
rect 41972 9998 42024 10004
rect 42156 10056 42208 10062
rect 42156 9998 42208 10004
rect 43076 10056 43128 10062
rect 43076 9998 43128 10004
rect 41236 9648 41288 9654
rect 41236 9590 41288 9596
rect 41340 9586 41368 9998
rect 41420 9920 41472 9926
rect 41420 9862 41472 9868
rect 41512 9920 41564 9926
rect 41512 9862 41564 9868
rect 40960 9580 41012 9586
rect 40960 9522 41012 9528
rect 41144 9580 41196 9586
rect 41144 9522 41196 9528
rect 41328 9580 41380 9586
rect 41328 9522 41380 9528
rect 39396 8628 39448 8634
rect 40144 8622 40356 8650
rect 39396 8570 39448 8576
rect 40040 8560 40092 8566
rect 40038 8528 40040 8537
rect 40092 8528 40094 8537
rect 39304 8492 39356 8498
rect 40038 8463 40094 8472
rect 40132 8492 40184 8498
rect 39304 8434 39356 8440
rect 40132 8434 40184 8440
rect 40224 8492 40276 8498
rect 40224 8434 40276 8440
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 38488 8266 38700 8294
rect 38384 7880 38436 7886
rect 38384 7822 38436 7828
rect 38396 7410 38424 7822
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 38396 6798 38424 7346
rect 38488 6866 38516 8266
rect 39132 7954 39160 8366
rect 40144 8362 40172 8434
rect 40040 8356 40092 8362
rect 40040 8298 40092 8304
rect 40132 8356 40184 8362
rect 40132 8298 40184 8304
rect 40052 7954 40080 8298
rect 39120 7948 39172 7954
rect 39120 7890 39172 7896
rect 40040 7948 40092 7954
rect 40040 7890 40092 7896
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 38384 6792 38436 6798
rect 38384 6734 38436 6740
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 38292 6656 38344 6662
rect 38290 6624 38292 6633
rect 38344 6624 38346 6633
rect 38290 6559 38346 6568
rect 40144 6390 40172 6734
rect 40236 6662 40264 8434
rect 40224 6656 40276 6662
rect 40224 6598 40276 6604
rect 38568 6384 38620 6390
rect 40132 6384 40184 6390
rect 38620 6332 38700 6338
rect 38568 6326 38700 6332
rect 40132 6326 40184 6332
rect 38580 6310 38700 6326
rect 38566 6216 38622 6225
rect 38566 6151 38568 6160
rect 38620 6151 38622 6160
rect 38568 6122 38620 6128
rect 38200 5704 38252 5710
rect 38200 5646 38252 5652
rect 37924 5160 37976 5166
rect 37924 5102 37976 5108
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37936 2990 37964 5102
rect 38212 3534 38240 5646
rect 38672 4826 38700 6310
rect 39396 6316 39448 6322
rect 39396 6258 39448 6264
rect 39408 6225 39436 6258
rect 39394 6216 39450 6225
rect 39394 6151 39396 6160
rect 39448 6151 39450 6160
rect 39396 6122 39448 6128
rect 39212 6112 39264 6118
rect 39408 6091 39436 6122
rect 39212 6054 39264 6060
rect 39224 5302 39252 6054
rect 40224 5636 40276 5642
rect 40224 5578 40276 5584
rect 40236 5302 40264 5578
rect 40328 5370 40356 8622
rect 40868 8628 40920 8634
rect 40868 8570 40920 8576
rect 40776 8560 40828 8566
rect 40776 8502 40828 8508
rect 40500 8492 40552 8498
rect 40500 8434 40552 8440
rect 40512 8378 40540 8434
rect 40512 8350 40632 8378
rect 40604 8090 40632 8350
rect 40592 8084 40644 8090
rect 40592 8026 40644 8032
rect 40408 6792 40460 6798
rect 40408 6734 40460 6740
rect 40420 6458 40448 6734
rect 40408 6452 40460 6458
rect 40408 6394 40460 6400
rect 40604 6338 40632 8026
rect 40684 7948 40736 7954
rect 40684 7890 40736 7896
rect 40696 7478 40724 7890
rect 40684 7472 40736 7478
rect 40684 7414 40736 7420
rect 40788 6644 40816 8502
rect 40880 8362 40908 8570
rect 40972 8401 41000 9522
rect 41156 8634 41184 9522
rect 41340 9382 41368 9522
rect 41328 9376 41380 9382
rect 41328 9318 41380 9324
rect 41432 9178 41460 9862
rect 41524 9586 41552 9862
rect 41512 9580 41564 9586
rect 41512 9522 41564 9528
rect 41984 9518 42012 9998
rect 42168 9722 42196 9998
rect 42156 9716 42208 9722
rect 42156 9658 42208 9664
rect 41972 9512 42024 9518
rect 41972 9454 42024 9460
rect 41420 9172 41472 9178
rect 41420 9114 41472 9120
rect 42156 9104 42208 9110
rect 42156 9046 42208 9052
rect 42168 8838 42196 9046
rect 42524 9036 42576 9042
rect 42524 8978 42576 8984
rect 42156 8832 42208 8838
rect 42156 8774 42208 8780
rect 41144 8628 41196 8634
rect 41144 8570 41196 8576
rect 42536 8566 42564 8978
rect 42616 8832 42668 8838
rect 42616 8774 42668 8780
rect 42524 8560 42576 8566
rect 42524 8502 42576 8508
rect 42248 8424 42300 8430
rect 40958 8392 41014 8401
rect 40868 8356 40920 8362
rect 42248 8366 42300 8372
rect 40958 8327 41014 8336
rect 41420 8356 41472 8362
rect 40868 8298 40920 8304
rect 40972 6798 41000 8327
rect 41420 8298 41472 8304
rect 40960 6792 41012 6798
rect 40960 6734 41012 6740
rect 41052 6724 41104 6730
rect 41052 6666 41104 6672
rect 40868 6656 40920 6662
rect 40788 6616 40868 6644
rect 40868 6598 40920 6604
rect 40960 6656 41012 6662
rect 40960 6598 41012 6604
rect 40420 6310 40632 6338
rect 40420 5642 40448 6310
rect 40880 6254 40908 6598
rect 40868 6248 40920 6254
rect 40868 6190 40920 6196
rect 40408 5636 40460 5642
rect 40408 5578 40460 5584
rect 40868 5636 40920 5642
rect 40868 5578 40920 5584
rect 40316 5364 40368 5370
rect 40316 5306 40368 5312
rect 39212 5296 39264 5302
rect 39212 5238 39264 5244
rect 40224 5296 40276 5302
rect 40224 5238 40276 5244
rect 40132 5024 40184 5030
rect 40132 4966 40184 4972
rect 38660 4820 38712 4826
rect 38660 4762 38712 4768
rect 39776 4690 40080 4706
rect 39764 4684 40092 4690
rect 39816 4678 40040 4684
rect 39764 4626 39816 4632
rect 40040 4626 40092 4632
rect 40144 4622 40172 4966
rect 40316 4752 40368 4758
rect 40316 4694 40368 4700
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 40132 4616 40184 4622
rect 40132 4558 40184 4564
rect 38566 4176 38622 4185
rect 38384 4140 38436 4146
rect 38566 4111 38568 4120
rect 38384 4082 38436 4088
rect 38620 4111 38622 4120
rect 38752 4140 38804 4146
rect 38568 4082 38620 4088
rect 38752 4082 38804 4088
rect 38396 3738 38424 4082
rect 38764 4010 38792 4082
rect 38752 4004 38804 4010
rect 38752 3946 38804 3952
rect 38844 3936 38896 3942
rect 38844 3878 38896 3884
rect 38384 3732 38436 3738
rect 38384 3674 38436 3680
rect 38200 3528 38252 3534
rect 38120 3488 38200 3516
rect 38120 3058 38148 3488
rect 38200 3470 38252 3476
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 38304 3058 38332 3470
rect 38856 3126 38884 3878
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39408 3194 39436 3674
rect 39868 3466 39896 4558
rect 40144 3534 40172 4558
rect 40328 4554 40356 4694
rect 40776 4684 40828 4690
rect 40776 4626 40828 4632
rect 40316 4548 40368 4554
rect 40316 4490 40368 4496
rect 40788 4214 40816 4626
rect 40776 4208 40828 4214
rect 40880 4185 40908 5578
rect 40972 5574 41000 6598
rect 40960 5568 41012 5574
rect 40960 5510 41012 5516
rect 41064 5302 41092 6666
rect 41234 5808 41290 5817
rect 41234 5743 41290 5752
rect 41248 5710 41276 5743
rect 41236 5704 41288 5710
rect 41236 5646 41288 5652
rect 41432 5556 41460 8298
rect 42260 8090 42288 8366
rect 42248 8084 42300 8090
rect 42248 8026 42300 8032
rect 42628 7818 42656 8774
rect 42800 8492 42852 8498
rect 42800 8434 42852 8440
rect 42708 7948 42760 7954
rect 42708 7890 42760 7896
rect 42616 7812 42668 7818
rect 42616 7754 42668 7760
rect 42720 7274 42748 7890
rect 42812 7750 42840 8434
rect 42800 7744 42852 7750
rect 42800 7686 42852 7692
rect 42708 7268 42760 7274
rect 42708 7210 42760 7216
rect 41880 6928 41932 6934
rect 41880 6870 41932 6876
rect 41696 6792 41748 6798
rect 41616 6752 41696 6780
rect 41616 6254 41644 6752
rect 41696 6734 41748 6740
rect 41694 6624 41750 6633
rect 41694 6559 41750 6568
rect 41604 6248 41656 6254
rect 41604 6190 41656 6196
rect 41708 6118 41736 6559
rect 41892 6322 41920 6870
rect 42720 6848 42748 7210
rect 42996 6866 43208 6882
rect 42892 6860 42944 6866
rect 42720 6820 42892 6848
rect 41972 6792 42024 6798
rect 41972 6734 42024 6740
rect 41880 6316 41932 6322
rect 41880 6258 41932 6264
rect 41512 6112 41564 6118
rect 41512 6054 41564 6060
rect 41696 6112 41748 6118
rect 41696 6054 41748 6060
rect 41524 5710 41552 6054
rect 41984 5930 42012 6734
rect 42720 6186 42748 6820
rect 42892 6802 42944 6808
rect 42996 6860 43220 6866
rect 42996 6854 43168 6860
rect 42996 6798 43024 6854
rect 43168 6802 43220 6808
rect 42984 6792 43036 6798
rect 42984 6734 43036 6740
rect 43076 6792 43128 6798
rect 43076 6734 43128 6740
rect 43088 6322 43116 6734
rect 43352 6724 43404 6730
rect 43352 6666 43404 6672
rect 43076 6316 43128 6322
rect 43076 6258 43128 6264
rect 43260 6248 43312 6254
rect 43260 6190 43312 6196
rect 42708 6180 42760 6186
rect 42708 6122 42760 6128
rect 41892 5914 42012 5930
rect 41880 5908 42012 5914
rect 41932 5902 42012 5908
rect 41880 5850 41932 5856
rect 43272 5778 43300 6190
rect 43364 5846 43392 6666
rect 43548 6322 43576 16546
rect 43720 16526 43772 16532
rect 43812 16584 43864 16590
rect 43812 16526 43864 16532
rect 43732 16114 43760 16526
rect 43824 16182 43852 16526
rect 43812 16176 43864 16182
rect 43812 16118 43864 16124
rect 43720 16108 43772 16114
rect 43720 16050 43772 16056
rect 44008 15502 44036 16594
rect 45020 16522 45048 16594
rect 45480 16522 45508 16594
rect 46572 16584 46624 16590
rect 46572 16526 46624 16532
rect 45008 16516 45060 16522
rect 45008 16458 45060 16464
rect 45100 16516 45152 16522
rect 45100 16458 45152 16464
rect 45468 16516 45520 16522
rect 45468 16458 45520 16464
rect 45112 15910 45140 16458
rect 45284 16448 45336 16454
rect 45284 16390 45336 16396
rect 45296 16250 45324 16390
rect 45284 16244 45336 16250
rect 45284 16186 45336 16192
rect 45192 16108 45244 16114
rect 45192 16050 45244 16056
rect 45204 15910 45232 16050
rect 46584 15978 46612 16526
rect 47032 16516 47084 16522
rect 47032 16458 47084 16464
rect 47044 16250 47072 16458
rect 47032 16244 47084 16250
rect 47032 16186 47084 16192
rect 46940 16108 46992 16114
rect 46940 16050 46992 16056
rect 46952 15994 46980 16050
rect 46572 15972 46624 15978
rect 46952 15966 47072 15994
rect 46572 15914 46624 15920
rect 45100 15904 45152 15910
rect 45100 15846 45152 15852
rect 45192 15904 45244 15910
rect 45192 15846 45244 15852
rect 43996 15496 44048 15502
rect 43996 15438 44048 15444
rect 43720 15088 43772 15094
rect 43720 15030 43772 15036
rect 43732 14550 43760 15030
rect 44008 15026 44036 15438
rect 44364 15360 44416 15366
rect 44364 15302 44416 15308
rect 46940 15360 46992 15366
rect 46940 15302 46992 15308
rect 44376 15026 44404 15302
rect 46952 15094 46980 15302
rect 47044 15162 47072 15966
rect 47136 15910 47164 17478
rect 47584 16108 47636 16114
rect 47584 16050 47636 16056
rect 47124 15904 47176 15910
rect 47124 15846 47176 15852
rect 47136 15502 47164 15846
rect 47596 15570 47624 16050
rect 47584 15564 47636 15570
rect 47584 15506 47636 15512
rect 47124 15496 47176 15502
rect 47124 15438 47176 15444
rect 47032 15156 47084 15162
rect 47032 15098 47084 15104
rect 46940 15088 46992 15094
rect 46940 15030 46992 15036
rect 43996 15020 44048 15026
rect 43996 14962 44048 14968
rect 44364 15020 44416 15026
rect 44364 14962 44416 14968
rect 46664 15020 46716 15026
rect 46664 14962 46716 14968
rect 44180 14816 44232 14822
rect 44180 14758 44232 14764
rect 43720 14544 43772 14550
rect 43720 14486 43772 14492
rect 44088 13524 44140 13530
rect 44088 13466 44140 13472
rect 44100 12850 44128 13466
rect 44192 13394 44220 14758
rect 44456 14408 44508 14414
rect 44456 14350 44508 14356
rect 44468 14006 44496 14350
rect 46296 14340 46348 14346
rect 46296 14282 46348 14288
rect 44456 14000 44508 14006
rect 44456 13942 44508 13948
rect 44364 13864 44416 13870
rect 44364 13806 44416 13812
rect 44180 13388 44232 13394
rect 44180 13330 44232 13336
rect 44192 12850 44220 13330
rect 44376 13326 44404 13806
rect 44468 13530 44496 13942
rect 45008 13932 45060 13938
rect 45008 13874 45060 13880
rect 44456 13524 44508 13530
rect 44456 13466 44508 13472
rect 44364 13320 44416 13326
rect 44364 13262 44416 13268
rect 44088 12844 44140 12850
rect 44088 12786 44140 12792
rect 44180 12844 44232 12850
rect 44180 12786 44232 12792
rect 44100 12209 44128 12786
rect 44192 12374 44220 12786
rect 44272 12708 44324 12714
rect 44272 12650 44324 12656
rect 44284 12442 44312 12650
rect 44272 12436 44324 12442
rect 44272 12378 44324 12384
rect 44180 12368 44232 12374
rect 44180 12310 44232 12316
rect 44086 12200 44142 12209
rect 44284 12170 44312 12378
rect 44086 12135 44142 12144
rect 44272 12164 44324 12170
rect 43720 12096 43772 12102
rect 43720 12038 43772 12044
rect 43732 11150 43760 12038
rect 44100 11626 44128 12135
rect 44272 12106 44324 12112
rect 44376 12102 44404 13262
rect 44640 13252 44692 13258
rect 44640 13194 44692 13200
rect 44652 12918 44680 13194
rect 44640 12912 44692 12918
rect 44640 12854 44692 12860
rect 45020 12434 45048 13874
rect 45468 13728 45520 13734
rect 45468 13670 45520 13676
rect 46204 13728 46256 13734
rect 46204 13670 46256 13676
rect 45480 13462 45508 13670
rect 45468 13456 45520 13462
rect 45468 13398 45520 13404
rect 44836 12406 45048 12434
rect 44364 12096 44416 12102
rect 44364 12038 44416 12044
rect 44836 11830 44864 12406
rect 44916 12232 44968 12238
rect 44916 12174 44968 12180
rect 44824 11824 44876 11830
rect 44824 11766 44876 11772
rect 44088 11620 44140 11626
rect 44088 11562 44140 11568
rect 43720 11144 43772 11150
rect 43720 11086 43772 11092
rect 44548 10804 44600 10810
rect 44548 10746 44600 10752
rect 43904 9920 43956 9926
rect 43904 9862 43956 9868
rect 43720 8492 43772 8498
rect 43720 8434 43772 8440
rect 43732 7410 43760 8434
rect 43812 8356 43864 8362
rect 43812 8298 43864 8304
rect 43720 7404 43772 7410
rect 43720 7346 43772 7352
rect 43732 6730 43760 7346
rect 43720 6724 43772 6730
rect 43720 6666 43772 6672
rect 43536 6316 43588 6322
rect 43536 6258 43588 6264
rect 43732 6254 43760 6666
rect 43720 6248 43772 6254
rect 43720 6190 43772 6196
rect 43352 5840 43404 5846
rect 43350 5808 43352 5817
rect 43404 5808 43406 5817
rect 43260 5772 43312 5778
rect 43350 5743 43406 5752
rect 43260 5714 43312 5720
rect 41512 5704 41564 5710
rect 41512 5646 41564 5652
rect 41972 5704 42024 5710
rect 41972 5646 42024 5652
rect 41984 5574 42012 5646
rect 43732 5574 43760 6190
rect 41972 5568 42024 5574
rect 41432 5528 41552 5556
rect 41052 5296 41104 5302
rect 41052 5238 41104 5244
rect 41064 4282 41092 5238
rect 41236 4480 41288 4486
rect 41236 4422 41288 4428
rect 41052 4276 41104 4282
rect 41052 4218 41104 4224
rect 40776 4150 40828 4156
rect 40866 4176 40922 4185
rect 41248 4146 41276 4422
rect 40866 4111 40922 4120
rect 41052 4140 41104 4146
rect 40880 4010 40908 4111
rect 41052 4082 41104 4088
rect 41236 4140 41288 4146
rect 41236 4082 41288 4088
rect 40868 4004 40920 4010
rect 40868 3946 40920 3952
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40776 3528 40828 3534
rect 40776 3470 40828 3476
rect 39856 3460 39908 3466
rect 39856 3402 39908 3408
rect 39580 3392 39632 3398
rect 39580 3334 39632 3340
rect 39672 3392 39724 3398
rect 39672 3334 39724 3340
rect 39592 3233 39620 3334
rect 39578 3224 39634 3233
rect 39396 3188 39448 3194
rect 39578 3159 39634 3168
rect 39396 3130 39448 3136
rect 38844 3120 38896 3126
rect 38844 3062 38896 3068
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 37924 2984 37976 2990
rect 37922 2952 37924 2961
rect 37976 2952 37978 2961
rect 37922 2887 37978 2896
rect 38200 2848 38252 2854
rect 38200 2790 38252 2796
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37648 1556 37700 1562
rect 37648 1498 37700 1504
rect 37752 800 37780 2314
rect 37832 2304 37884 2310
rect 37832 2246 37884 2252
rect 37844 2038 37872 2246
rect 37832 2032 37884 2038
rect 37832 1974 37884 1980
rect 38212 800 38240 2790
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 38752 2304 38804 2310
rect 38752 2246 38804 2252
rect 38764 1494 38792 2246
rect 38752 1488 38804 1494
rect 38752 1430 38804 1436
rect 39224 800 39252 2314
rect 39684 800 39712 3334
rect 39868 3194 39896 3402
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39868 3058 39896 3130
rect 40788 3058 40816 3470
rect 40880 3398 40908 3946
rect 40960 3936 41012 3942
rect 40960 3878 41012 3884
rect 40868 3392 40920 3398
rect 40868 3334 40920 3340
rect 40866 3224 40922 3233
rect 40866 3159 40922 3168
rect 40880 3058 40908 3159
rect 39856 3052 39908 3058
rect 39856 2994 39908 3000
rect 40776 3052 40828 3058
rect 40776 2994 40828 3000
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 40972 2774 41000 3878
rect 41064 3126 41092 4082
rect 41248 3534 41276 4082
rect 41328 4004 41380 4010
rect 41328 3946 41380 3952
rect 41420 4004 41472 4010
rect 41420 3946 41472 3952
rect 41340 3777 41368 3946
rect 41326 3768 41382 3777
rect 41432 3738 41460 3946
rect 41326 3703 41382 3712
rect 41420 3732 41472 3738
rect 41420 3674 41472 3680
rect 41524 3534 41552 5528
rect 41972 5510 42024 5516
rect 43720 5568 43772 5574
rect 43720 5510 43772 5516
rect 41984 5098 42012 5510
rect 41972 5092 42024 5098
rect 41972 5034 42024 5040
rect 41984 4078 42012 5034
rect 43824 4282 43852 8298
rect 43916 7750 43944 9862
rect 43904 7744 43956 7750
rect 43904 7686 43956 7692
rect 43812 4276 43864 4282
rect 43812 4218 43864 4224
rect 41972 4072 42024 4078
rect 41972 4014 42024 4020
rect 42432 4072 42484 4078
rect 42432 4014 42484 4020
rect 42154 3632 42210 3641
rect 42154 3567 42156 3576
rect 42208 3567 42210 3576
rect 42156 3538 42208 3544
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 41512 3528 41564 3534
rect 41512 3470 41564 3476
rect 42248 3528 42300 3534
rect 42248 3470 42300 3476
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 41340 3194 41368 3402
rect 41788 3392 41840 3398
rect 41788 3334 41840 3340
rect 41328 3188 41380 3194
rect 41328 3130 41380 3136
rect 41800 3126 41828 3334
rect 42260 3194 42288 3470
rect 42248 3188 42300 3194
rect 42248 3130 42300 3136
rect 41052 3120 41104 3126
rect 41052 3062 41104 3068
rect 41788 3120 41840 3126
rect 41788 3062 41840 3068
rect 41144 3052 41196 3058
rect 41144 2994 41196 3000
rect 41156 2922 41184 2994
rect 42444 2990 42472 4014
rect 42798 3768 42854 3777
rect 42798 3703 42800 3712
rect 42852 3703 42854 3712
rect 43442 3768 43498 3777
rect 43442 3703 43498 3712
rect 42800 3674 42852 3680
rect 43456 3670 43484 3703
rect 43444 3664 43496 3670
rect 42536 3590 42840 3618
rect 43444 3606 43496 3612
rect 42536 3534 42564 3590
rect 42812 3534 42840 3590
rect 43824 3534 43852 4218
rect 42524 3528 42576 3534
rect 42708 3528 42760 3534
rect 42524 3470 42576 3476
rect 42628 3488 42708 3516
rect 42432 2984 42484 2990
rect 42432 2926 42484 2932
rect 41144 2916 41196 2922
rect 41144 2858 41196 2864
rect 42628 2854 42656 3488
rect 42708 3470 42760 3476
rect 42800 3528 42852 3534
rect 42800 3470 42852 3476
rect 43812 3528 43864 3534
rect 43812 3470 43864 3476
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42720 3233 42748 3334
rect 42706 3224 42762 3233
rect 42706 3159 42762 3168
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 40972 2746 41184 2774
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40604 800 40632 2314
rect 41156 800 41184 2746
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 2106 41368 2450
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 41328 2100 41380 2106
rect 41328 2042 41380 2048
rect 42076 800 42104 2314
rect 42628 870 42748 898
rect 42628 800 42656 870
rect 20272 734 20576 762
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 42720 762 42748 870
rect 42996 762 43024 3334
rect 43916 3058 43944 7686
rect 44560 7410 44588 10746
rect 44548 7404 44600 7410
rect 44548 7346 44600 7352
rect 44836 5692 44864 11766
rect 44928 11558 44956 12174
rect 44916 11552 44968 11558
rect 44916 11494 44968 11500
rect 45480 9654 45508 13398
rect 46216 13326 46244 13670
rect 46308 13530 46336 14282
rect 46676 14074 46704 14962
rect 46664 14068 46716 14074
rect 46664 14010 46716 14016
rect 46296 13524 46348 13530
rect 46296 13466 46348 13472
rect 46204 13320 46256 13326
rect 46204 13262 46256 13268
rect 45652 12844 45704 12850
rect 45652 12786 45704 12792
rect 45560 12640 45612 12646
rect 45560 12582 45612 12588
rect 45572 12238 45600 12582
rect 45560 12232 45612 12238
rect 45560 12174 45612 12180
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45572 11082 45600 12038
rect 45664 11626 45692 12786
rect 46676 12714 46704 14010
rect 47872 12918 47900 17546
rect 47952 16448 48004 16454
rect 47952 16390 48004 16396
rect 47964 16182 47992 16390
rect 47952 16176 48004 16182
rect 47952 16118 48004 16124
rect 48412 16108 48464 16114
rect 48412 16050 48464 16056
rect 47952 15428 48004 15434
rect 47952 15370 48004 15376
rect 47964 15026 47992 15370
rect 47952 15020 48004 15026
rect 47952 14962 48004 14968
rect 47964 14278 47992 14962
rect 48424 14414 48452 16050
rect 48412 14408 48464 14414
rect 48412 14350 48464 14356
rect 47952 14272 48004 14278
rect 47952 14214 48004 14220
rect 47964 13870 47992 14214
rect 47952 13864 48004 13870
rect 47952 13806 48004 13812
rect 48044 13456 48096 13462
rect 48044 13398 48096 13404
rect 48056 12986 48084 13398
rect 48044 12980 48096 12986
rect 48044 12922 48096 12928
rect 47860 12912 47912 12918
rect 47860 12854 47912 12860
rect 48228 12912 48280 12918
rect 48228 12854 48280 12860
rect 45744 12708 45796 12714
rect 45744 12650 45796 12656
rect 46664 12708 46716 12714
rect 46664 12650 46716 12656
rect 45756 11830 45784 12650
rect 45744 11824 45796 11830
rect 45744 11766 45796 11772
rect 45652 11620 45704 11626
rect 45652 11562 45704 11568
rect 48240 11558 48268 12854
rect 48424 12782 48452 14350
rect 48412 12776 48464 12782
rect 48412 12718 48464 12724
rect 48424 12434 48452 12718
rect 48332 12406 48452 12434
rect 48228 11552 48280 11558
rect 48228 11494 48280 11500
rect 47676 11348 47728 11354
rect 47676 11290 47728 11296
rect 45560 11076 45612 11082
rect 45560 11018 45612 11024
rect 45572 10130 45600 11018
rect 47688 10266 47716 11290
rect 48332 11082 48360 12406
rect 48608 12306 48636 17818
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 54772 15706 54800 39374
rect 54760 15700 54812 15706
rect 54760 15642 54812 15648
rect 53104 15496 53156 15502
rect 53104 15438 53156 15444
rect 53012 15428 53064 15434
rect 53012 15370 53064 15376
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 53024 15162 53052 15370
rect 53012 15156 53064 15162
rect 53012 15098 53064 15104
rect 50620 14340 50672 14346
rect 50620 14282 50672 14288
rect 50160 14272 50212 14278
rect 50160 14214 50212 14220
rect 50172 13326 50200 14214
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 50632 14074 50660 14282
rect 50620 14068 50672 14074
rect 50620 14010 50672 14016
rect 50528 13932 50580 13938
rect 50528 13874 50580 13880
rect 50620 13932 50672 13938
rect 50620 13874 50672 13880
rect 50540 13530 50568 13874
rect 50528 13524 50580 13530
rect 50528 13466 50580 13472
rect 49148 13320 49200 13326
rect 49148 13262 49200 13268
rect 50160 13320 50212 13326
rect 50160 13262 50212 13268
rect 49160 12442 49188 13262
rect 49240 13184 49292 13190
rect 49240 13126 49292 13132
rect 49252 12918 49280 13126
rect 49240 12912 49292 12918
rect 49240 12854 49292 12860
rect 49148 12436 49200 12442
rect 49148 12378 49200 12384
rect 48596 12300 48648 12306
rect 48596 12242 48648 12248
rect 49700 12232 49752 12238
rect 49700 12174 49752 12180
rect 49712 12102 49740 12174
rect 50172 12170 50200 13262
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50632 12442 50660 13874
rect 53116 13870 53144 15438
rect 53196 15020 53248 15026
rect 53196 14962 53248 14968
rect 53208 14006 53236 14962
rect 54024 14408 54076 14414
rect 54024 14350 54076 14356
rect 53748 14272 53800 14278
rect 53748 14214 53800 14220
rect 53760 14006 53788 14214
rect 53196 14000 53248 14006
rect 53196 13942 53248 13948
rect 53748 14000 53800 14006
rect 53748 13942 53800 13948
rect 52644 13864 52696 13870
rect 52644 13806 52696 13812
rect 53104 13864 53156 13870
rect 53104 13806 53156 13812
rect 50988 13320 51040 13326
rect 50988 13262 51040 13268
rect 51000 12986 51028 13262
rect 52656 12986 52684 13806
rect 53748 13320 53800 13326
rect 53748 13262 53800 13268
rect 50988 12980 51040 12986
rect 50988 12922 51040 12928
rect 52644 12980 52696 12986
rect 52644 12922 52696 12928
rect 50804 12844 50856 12850
rect 50804 12786 50856 12792
rect 50620 12436 50672 12442
rect 50620 12378 50672 12384
rect 50160 12164 50212 12170
rect 50160 12106 50212 12112
rect 50816 12102 50844 12786
rect 50896 12776 50948 12782
rect 50896 12718 50948 12724
rect 50908 12374 50936 12718
rect 50896 12368 50948 12374
rect 50896 12310 50948 12316
rect 49700 12096 49752 12102
rect 49700 12038 49752 12044
rect 50804 12096 50856 12102
rect 50804 12038 50856 12044
rect 48504 11824 48556 11830
rect 48504 11766 48556 11772
rect 48320 11076 48372 11082
rect 48320 11018 48372 11024
rect 48516 10810 48544 11766
rect 49712 11762 49740 12038
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 49700 11756 49752 11762
rect 49700 11698 49752 11704
rect 48596 11552 48648 11558
rect 48596 11494 48648 11500
rect 48608 11354 48636 11494
rect 48596 11348 48648 11354
rect 48596 11290 48648 11296
rect 49884 11008 49936 11014
rect 49884 10950 49936 10956
rect 48504 10804 48556 10810
rect 48504 10746 48556 10752
rect 49896 10742 49924 10950
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 50816 10810 50844 12038
rect 50908 11354 50936 12310
rect 50988 12096 51040 12102
rect 50988 12038 51040 12044
rect 52000 12096 52052 12102
rect 52000 12038 52052 12044
rect 50896 11348 50948 11354
rect 50896 11290 50948 11296
rect 50804 10804 50856 10810
rect 50804 10746 50856 10752
rect 48596 10736 48648 10742
rect 48596 10678 48648 10684
rect 49884 10736 49936 10742
rect 49884 10678 49936 10684
rect 49976 10736 50028 10742
rect 49976 10678 50028 10684
rect 48228 10600 48280 10606
rect 48228 10542 48280 10548
rect 47676 10260 47728 10266
rect 47676 10202 47728 10208
rect 45560 10124 45612 10130
rect 45612 10084 45692 10112
rect 45560 10066 45612 10072
rect 45560 9988 45612 9994
rect 45560 9930 45612 9936
rect 45468 9648 45520 9654
rect 45468 9590 45520 9596
rect 45572 9450 45600 9930
rect 45560 9444 45612 9450
rect 45560 9386 45612 9392
rect 45192 9376 45244 9382
rect 45192 9318 45244 9324
rect 45204 8974 45232 9318
rect 45192 8968 45244 8974
rect 45192 8910 45244 8916
rect 45008 8832 45060 8838
rect 45008 8774 45060 8780
rect 45020 8566 45048 8774
rect 45008 8560 45060 8566
rect 45664 8514 45692 10084
rect 47032 9920 47084 9926
rect 47032 9862 47084 9868
rect 47044 9586 47072 9862
rect 48240 9586 48268 10542
rect 47032 9580 47084 9586
rect 47032 9522 47084 9528
rect 48228 9580 48280 9586
rect 48228 9522 48280 9528
rect 46940 9104 46992 9110
rect 46940 9046 46992 9052
rect 45008 8502 45060 8508
rect 45572 8498 45692 8514
rect 45560 8492 45692 8498
rect 45612 8486 45692 8492
rect 45560 8434 45612 8440
rect 46952 8362 46980 9046
rect 47044 9042 47072 9522
rect 48608 9518 48636 10678
rect 49608 10260 49660 10266
rect 49608 10202 49660 10208
rect 49620 9518 49648 10202
rect 49988 9586 50016 10678
rect 51000 10470 51028 12038
rect 51540 11824 51592 11830
rect 51540 11766 51592 11772
rect 51552 11354 51580 11766
rect 52012 11626 52040 12038
rect 52000 11620 52052 11626
rect 52000 11562 52052 11568
rect 51816 11552 51868 11558
rect 51816 11494 51868 11500
rect 51540 11348 51592 11354
rect 51540 11290 51592 11296
rect 50068 10464 50120 10470
rect 50068 10406 50120 10412
rect 50988 10464 51040 10470
rect 50988 10406 51040 10412
rect 49976 9580 50028 9586
rect 49976 9522 50028 9528
rect 48596 9512 48648 9518
rect 48596 9454 48648 9460
rect 49516 9512 49568 9518
rect 49516 9454 49568 9460
rect 49608 9512 49660 9518
rect 49608 9454 49660 9460
rect 47032 9036 47084 9042
rect 47032 8978 47084 8984
rect 46940 8356 46992 8362
rect 46940 8298 46992 8304
rect 47768 8356 47820 8362
rect 47768 8298 47820 8304
rect 45192 7812 45244 7818
rect 45192 7754 45244 7760
rect 45204 7206 45232 7754
rect 45284 7404 45336 7410
rect 45284 7346 45336 7352
rect 47308 7404 47360 7410
rect 47308 7346 47360 7352
rect 45192 7200 45244 7206
rect 45192 7142 45244 7148
rect 45100 5704 45152 5710
rect 44836 5664 45100 5692
rect 45100 5646 45152 5652
rect 45112 4554 45140 5646
rect 45100 4548 45152 4554
rect 45100 4490 45152 4496
rect 45204 3534 45232 7142
rect 45296 5574 45324 7346
rect 46940 7336 46992 7342
rect 46940 7278 46992 7284
rect 46204 7200 46256 7206
rect 46204 7142 46256 7148
rect 46572 7200 46624 7206
rect 46572 7142 46624 7148
rect 45560 6792 45612 6798
rect 45560 6734 45612 6740
rect 45572 6118 45600 6734
rect 46216 6730 46244 7142
rect 46584 7002 46612 7142
rect 46572 6996 46624 7002
rect 46572 6938 46624 6944
rect 46572 6792 46624 6798
rect 46624 6752 46888 6780
rect 46572 6734 46624 6740
rect 46204 6724 46256 6730
rect 46204 6666 46256 6672
rect 46572 6316 46624 6322
rect 46572 6258 46624 6264
rect 46664 6316 46716 6322
rect 46664 6258 46716 6264
rect 45560 6112 45612 6118
rect 45560 6054 45612 6060
rect 46584 5778 46612 6258
rect 46572 5772 46624 5778
rect 46572 5714 46624 5720
rect 46676 5710 46704 6258
rect 46860 6118 46888 6752
rect 46952 6458 46980 7278
rect 46940 6452 46992 6458
rect 46940 6394 46992 6400
rect 47032 6452 47084 6458
rect 47032 6394 47084 6400
rect 46756 6112 46808 6118
rect 46756 6054 46808 6060
rect 46848 6112 46900 6118
rect 46848 6054 46900 6060
rect 46664 5704 46716 5710
rect 46664 5646 46716 5652
rect 45652 5636 45704 5642
rect 45652 5578 45704 5584
rect 45284 5568 45336 5574
rect 45284 5510 45336 5516
rect 45468 4684 45520 4690
rect 45468 4626 45520 4632
rect 45480 4282 45508 4626
rect 45468 4276 45520 4282
rect 45468 4218 45520 4224
rect 45480 4146 45508 4218
rect 45468 4140 45520 4146
rect 45388 4100 45468 4128
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 43904 3052 43956 3058
rect 43904 2994 43956 3000
rect 44088 2848 44140 2854
rect 44088 2790 44140 2796
rect 43536 2372 43588 2378
rect 43536 2314 43588 2320
rect 43548 800 43576 2314
rect 44100 800 44128 2790
rect 45388 2446 45416 4100
rect 45468 4082 45520 4088
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45376 2440 45428 2446
rect 45376 2382 45428 2388
rect 45008 2304 45060 2310
rect 45008 2246 45060 2252
rect 45020 800 45048 2246
rect 45480 800 45508 3334
rect 45664 3058 45692 5578
rect 45742 5128 45798 5137
rect 45742 5063 45798 5072
rect 45756 4146 45784 5063
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 45834 4176 45890 4185
rect 45744 4140 45796 4146
rect 45834 4111 45836 4120
rect 45744 4082 45796 4088
rect 45888 4111 45890 4120
rect 45836 4082 45888 4088
rect 45652 3052 45704 3058
rect 45652 2994 45704 3000
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45664 2446 45692 2790
rect 45848 2446 45876 4082
rect 46308 3534 46336 4626
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46400 3670 46428 4150
rect 46388 3664 46440 3670
rect 46388 3606 46440 3612
rect 45928 3528 45980 3534
rect 45926 3496 45928 3505
rect 46296 3528 46348 3534
rect 45980 3496 45982 3505
rect 46296 3470 46348 3476
rect 45926 3431 45982 3440
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 46480 3392 46532 3398
rect 46480 3334 46532 3340
rect 45928 3052 45980 3058
rect 45928 2994 45980 3000
rect 45940 2650 45968 2994
rect 46492 2938 46520 3334
rect 46400 2910 46520 2938
rect 46400 2854 46428 2910
rect 46676 2854 46704 3402
rect 46768 2990 46796 6054
rect 47044 5846 47072 6394
rect 47320 6322 47348 7346
rect 47124 6316 47176 6322
rect 47124 6258 47176 6264
rect 47308 6316 47360 6322
rect 47308 6258 47360 6264
rect 47032 5840 47084 5846
rect 47032 5782 47084 5788
rect 47136 5778 47164 6258
rect 47490 6216 47546 6225
rect 47490 6151 47546 6160
rect 47504 5914 47532 6151
rect 47308 5908 47360 5914
rect 47492 5908 47544 5914
rect 47360 5868 47440 5896
rect 47308 5850 47360 5856
rect 47124 5772 47176 5778
rect 47124 5714 47176 5720
rect 47032 5636 47084 5642
rect 47032 5578 47084 5584
rect 47044 4214 47072 5578
rect 47136 4690 47164 5714
rect 47412 5710 47440 5868
rect 47492 5850 47544 5856
rect 47400 5704 47452 5710
rect 47400 5646 47452 5652
rect 47124 4684 47176 4690
rect 47124 4626 47176 4632
rect 47492 4684 47544 4690
rect 47492 4626 47544 4632
rect 47032 4208 47084 4214
rect 46846 4176 46902 4185
rect 47084 4168 47164 4196
rect 47032 4150 47084 4156
rect 46846 4111 46848 4120
rect 46900 4111 46902 4120
rect 46848 4082 46900 4088
rect 47032 3936 47084 3942
rect 47032 3878 47084 3884
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 46952 3398 46980 3470
rect 46940 3392 46992 3398
rect 46940 3334 46992 3340
rect 47044 3126 47072 3878
rect 47136 3534 47164 4168
rect 47504 3534 47532 4626
rect 47584 4140 47636 4146
rect 47584 4082 47636 4088
rect 47596 3942 47624 4082
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47582 3768 47638 3777
rect 47582 3703 47584 3712
rect 47636 3703 47638 3712
rect 47584 3674 47636 3680
rect 47582 3632 47638 3641
rect 47582 3567 47584 3576
rect 47636 3567 47638 3576
rect 47584 3538 47636 3544
rect 47124 3528 47176 3534
rect 47492 3528 47544 3534
rect 47124 3470 47176 3476
rect 47214 3496 47270 3505
rect 47492 3470 47544 3476
rect 47214 3431 47216 3440
rect 47268 3431 47270 3440
rect 47216 3402 47268 3408
rect 47032 3120 47084 3126
rect 47032 3062 47084 3068
rect 47780 3058 47808 8298
rect 49528 8022 49556 9454
rect 50080 8974 50108 10406
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50712 9716 50764 9722
rect 50712 9658 50764 9664
rect 50724 9178 50752 9658
rect 51828 9586 51856 11494
rect 52656 10606 52684 12922
rect 53760 12374 53788 13262
rect 54036 13190 54064 14350
rect 54576 14340 54628 14346
rect 54576 14282 54628 14288
rect 54116 13728 54168 13734
rect 54116 13670 54168 13676
rect 54128 13258 54156 13670
rect 54588 13530 54616 14282
rect 54576 13524 54628 13530
rect 54576 13466 54628 13472
rect 54944 13388 54996 13394
rect 54944 13330 54996 13336
rect 54116 13252 54168 13258
rect 54116 13194 54168 13200
rect 54024 13184 54076 13190
rect 54024 13126 54076 13132
rect 53840 12844 53892 12850
rect 53840 12786 53892 12792
rect 53852 12374 53880 12786
rect 54036 12782 54064 13126
rect 54024 12776 54076 12782
rect 54024 12718 54076 12724
rect 53932 12640 53984 12646
rect 53932 12582 53984 12588
rect 53748 12368 53800 12374
rect 53748 12310 53800 12316
rect 53840 12368 53892 12374
rect 53840 12310 53892 12316
rect 53760 12238 53788 12310
rect 53748 12232 53800 12238
rect 53748 12174 53800 12180
rect 53564 12096 53616 12102
rect 53564 12038 53616 12044
rect 53576 11898 53604 12038
rect 53564 11892 53616 11898
rect 53564 11834 53616 11840
rect 53656 11824 53708 11830
rect 53656 11766 53708 11772
rect 53104 11008 53156 11014
rect 53104 10950 53156 10956
rect 52644 10600 52696 10606
rect 52644 10542 52696 10548
rect 52656 9722 52684 10542
rect 52920 10124 52972 10130
rect 52920 10066 52972 10072
rect 52644 9716 52696 9722
rect 52644 9658 52696 9664
rect 51816 9580 51868 9586
rect 51816 9522 51868 9528
rect 50988 9512 51040 9518
rect 50988 9454 51040 9460
rect 50712 9172 50764 9178
rect 50712 9114 50764 9120
rect 50160 9104 50212 9110
rect 50160 9046 50212 9052
rect 50068 8968 50120 8974
rect 50068 8910 50120 8916
rect 50080 8634 50108 8910
rect 50068 8628 50120 8634
rect 50172 8616 50200 9046
rect 51000 8974 51028 9454
rect 50712 8968 50764 8974
rect 50712 8910 50764 8916
rect 50988 8968 51040 8974
rect 50988 8910 51040 8916
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50620 8628 50672 8634
rect 50172 8588 50292 8616
rect 50068 8570 50120 8576
rect 50160 8492 50212 8498
rect 50160 8434 50212 8440
rect 50172 8090 50200 8434
rect 50160 8084 50212 8090
rect 50160 8026 50212 8032
rect 49516 8016 49568 8022
rect 49516 7958 49568 7964
rect 50264 7886 50292 8588
rect 50620 8570 50672 8576
rect 50632 7954 50660 8570
rect 50724 8022 50752 8910
rect 52656 8566 52684 9658
rect 52932 8838 52960 10066
rect 53116 10062 53144 10950
rect 53288 10668 53340 10674
rect 53288 10610 53340 10616
rect 53300 10266 53328 10610
rect 53288 10260 53340 10266
rect 53288 10202 53340 10208
rect 53104 10056 53156 10062
rect 53104 9998 53156 10004
rect 53196 10056 53248 10062
rect 53196 9998 53248 10004
rect 53208 9654 53236 9998
rect 53564 9716 53616 9722
rect 53564 9658 53616 9664
rect 53196 9648 53248 9654
rect 53196 9590 53248 9596
rect 53576 9450 53604 9658
rect 53564 9444 53616 9450
rect 53564 9386 53616 9392
rect 53012 9376 53064 9382
rect 53012 9318 53064 9324
rect 53024 9178 53052 9318
rect 53012 9172 53064 9178
rect 53012 9114 53064 9120
rect 52920 8832 52972 8838
rect 52920 8774 52972 8780
rect 52644 8560 52696 8566
rect 52644 8502 52696 8508
rect 50712 8016 50764 8022
rect 50712 7958 50764 7964
rect 52656 7954 52684 8502
rect 50620 7948 50672 7954
rect 50620 7890 50672 7896
rect 52644 7948 52696 7954
rect 52644 7890 52696 7896
rect 50252 7880 50304 7886
rect 50252 7822 50304 7828
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 52932 7478 52960 8774
rect 53024 8430 53052 9114
rect 53288 8968 53340 8974
rect 53288 8910 53340 8916
rect 53300 8498 53328 8910
rect 53668 8906 53696 11766
rect 53944 11558 53972 12582
rect 54024 12232 54076 12238
rect 54024 12174 54076 12180
rect 54036 11762 54064 12174
rect 54128 12170 54156 13194
rect 54208 12844 54260 12850
rect 54208 12786 54260 12792
rect 54220 12238 54248 12786
rect 54956 12782 54984 13330
rect 55864 12980 55916 12986
rect 55864 12922 55916 12928
rect 55496 12912 55548 12918
rect 55496 12854 55548 12860
rect 55312 12844 55364 12850
rect 55312 12786 55364 12792
rect 54944 12776 54996 12782
rect 54944 12718 54996 12724
rect 54760 12640 54812 12646
rect 54760 12582 54812 12588
rect 55220 12640 55272 12646
rect 55220 12582 55272 12588
rect 54772 12238 54800 12582
rect 54208 12232 54260 12238
rect 54208 12174 54260 12180
rect 54760 12232 54812 12238
rect 54760 12174 54812 12180
rect 55232 12170 55260 12582
rect 55324 12442 55352 12786
rect 55312 12436 55364 12442
rect 55312 12378 55364 12384
rect 55508 12170 55536 12854
rect 55876 12782 55904 12922
rect 55864 12776 55916 12782
rect 55864 12718 55916 12724
rect 54116 12164 54168 12170
rect 54116 12106 54168 12112
rect 55220 12164 55272 12170
rect 55220 12106 55272 12112
rect 55496 12164 55548 12170
rect 55496 12106 55548 12112
rect 55876 11762 55904 12718
rect 54024 11756 54076 11762
rect 54024 11698 54076 11704
rect 55864 11756 55916 11762
rect 55864 11698 55916 11704
rect 53932 11552 53984 11558
rect 53932 11494 53984 11500
rect 53944 9994 53972 11494
rect 54392 11144 54444 11150
rect 54392 11086 54444 11092
rect 54404 10810 54432 11086
rect 54392 10804 54444 10810
rect 54392 10746 54444 10752
rect 53932 9988 53984 9994
rect 53932 9930 53984 9936
rect 54024 9580 54076 9586
rect 54024 9522 54076 9528
rect 53748 9376 53800 9382
rect 53748 9318 53800 9324
rect 53760 8906 53788 9318
rect 54036 9178 54064 9522
rect 54024 9172 54076 9178
rect 54024 9114 54076 9120
rect 53656 8900 53708 8906
rect 53656 8842 53708 8848
rect 53748 8900 53800 8906
rect 53748 8842 53800 8848
rect 53288 8492 53340 8498
rect 53288 8434 53340 8440
rect 53012 8424 53064 8430
rect 53012 8366 53064 8372
rect 53012 8288 53064 8294
rect 53012 8230 53064 8236
rect 52920 7472 52972 7478
rect 52920 7414 52972 7420
rect 53024 7410 53052 8230
rect 53300 8090 53328 8434
rect 53288 8084 53340 8090
rect 53288 8026 53340 8032
rect 53104 7812 53156 7818
rect 53104 7754 53156 7760
rect 53116 7546 53144 7754
rect 53104 7540 53156 7546
rect 53104 7482 53156 7488
rect 53012 7404 53064 7410
rect 53012 7346 53064 7352
rect 49148 6792 49200 6798
rect 49148 6734 49200 6740
rect 50620 6792 50672 6798
rect 50620 6734 50672 6740
rect 49160 6662 49188 6734
rect 49332 6724 49384 6730
rect 49332 6666 49384 6672
rect 47952 6656 48004 6662
rect 47952 6598 48004 6604
rect 49148 6656 49200 6662
rect 49148 6598 49200 6604
rect 47964 5574 47992 6598
rect 48872 6452 48924 6458
rect 48872 6394 48924 6400
rect 48044 6248 48096 6254
rect 48044 6190 48096 6196
rect 48056 5846 48084 6190
rect 48596 6112 48648 6118
rect 48596 6054 48648 6060
rect 48044 5840 48096 5846
rect 48044 5782 48096 5788
rect 47952 5568 48004 5574
rect 47952 5510 48004 5516
rect 47964 3670 47992 5510
rect 48608 5234 48636 6054
rect 48780 5636 48832 5642
rect 48780 5578 48832 5584
rect 48596 5228 48648 5234
rect 48596 5170 48648 5176
rect 48044 4684 48096 4690
rect 48044 4626 48096 4632
rect 48056 4146 48084 4626
rect 48320 4548 48372 4554
rect 48320 4490 48372 4496
rect 48044 4140 48096 4146
rect 48044 4082 48096 4088
rect 48044 4004 48096 4010
rect 48044 3946 48096 3952
rect 47952 3664 48004 3670
rect 47952 3606 48004 3612
rect 47860 3528 47912 3534
rect 47858 3496 47860 3505
rect 47912 3496 47914 3505
rect 48056 3466 48084 3946
rect 47858 3431 47914 3440
rect 48044 3460 48096 3466
rect 48044 3402 48096 3408
rect 48332 3398 48360 4490
rect 48502 3632 48558 3641
rect 48502 3567 48504 3576
rect 48556 3567 48558 3576
rect 48504 3538 48556 3544
rect 48320 3392 48372 3398
rect 48320 3334 48372 3340
rect 48412 3392 48464 3398
rect 48412 3334 48464 3340
rect 47768 3052 47820 3058
rect 47768 2994 47820 3000
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46940 2916 46992 2922
rect 46940 2858 46992 2864
rect 46388 2848 46440 2854
rect 46388 2790 46440 2796
rect 46664 2848 46716 2854
rect 46664 2790 46716 2796
rect 45928 2644 45980 2650
rect 45928 2586 45980 2592
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45744 2372 45796 2378
rect 45744 2314 45796 2320
rect 46756 2372 46808 2378
rect 46756 2314 46808 2320
rect 45756 1902 45784 2314
rect 45744 1896 45796 1902
rect 45744 1838 45796 1844
rect 46492 870 46612 898
rect 46492 800 46520 870
rect 42720 734 43024 762
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46584 762 46612 870
rect 46768 762 46796 2314
rect 46952 800 46980 2858
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 47964 800 47992 2382
rect 48228 2372 48280 2378
rect 48228 2314 48280 2320
rect 48136 2304 48188 2310
rect 48136 2246 48188 2252
rect 48148 2038 48176 2246
rect 48136 2032 48188 2038
rect 48136 1974 48188 1980
rect 48240 1698 48268 2314
rect 48228 1692 48280 1698
rect 48228 1634 48280 1640
rect 48424 800 48452 3334
rect 48608 3058 48636 5170
rect 48792 4826 48820 5578
rect 48884 5114 48912 6394
rect 49160 5710 49188 6598
rect 49148 5704 49200 5710
rect 49148 5646 49200 5652
rect 48884 5086 49096 5114
rect 48964 5024 49016 5030
rect 48964 4966 49016 4972
rect 48780 4820 48832 4826
rect 48780 4762 48832 4768
rect 48872 4752 48924 4758
rect 48872 4694 48924 4700
rect 48884 4622 48912 4694
rect 48688 4616 48740 4622
rect 48688 4558 48740 4564
rect 48872 4616 48924 4622
rect 48872 4558 48924 4564
rect 48700 4214 48728 4558
rect 48884 4282 48912 4558
rect 48976 4554 49004 4966
rect 48964 4548 49016 4554
rect 48964 4490 49016 4496
rect 48872 4276 48924 4282
rect 48872 4218 48924 4224
rect 48688 4208 48740 4214
rect 48688 4150 48740 4156
rect 48700 3194 48728 4150
rect 49068 4146 49096 5086
rect 49148 4616 49200 4622
rect 49148 4558 49200 4564
rect 49160 4146 49188 4558
rect 48780 4140 48832 4146
rect 48780 4082 48832 4088
rect 49056 4140 49108 4146
rect 49056 4082 49108 4088
rect 49148 4140 49200 4146
rect 49148 4082 49200 4088
rect 48688 3188 48740 3194
rect 48688 3130 48740 3136
rect 48596 3052 48648 3058
rect 48596 2994 48648 3000
rect 48792 2961 48820 4082
rect 48872 3528 48924 3534
rect 48870 3496 48872 3505
rect 48924 3496 48926 3505
rect 48870 3431 48926 3440
rect 48778 2952 48834 2961
rect 48778 2887 48834 2896
rect 48792 2854 48820 2887
rect 48780 2848 48832 2854
rect 48780 2790 48832 2796
rect 49068 2582 49096 4082
rect 49344 4010 49372 6666
rect 49424 6656 49476 6662
rect 49424 6598 49476 6604
rect 49436 6118 49464 6598
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 49424 6112 49476 6118
rect 49424 6054 49476 6060
rect 50160 6112 50212 6118
rect 50160 6054 50212 6060
rect 50172 5574 50200 6054
rect 50632 5914 50660 6734
rect 52644 6656 52696 6662
rect 52644 6598 52696 6604
rect 50620 5908 50672 5914
rect 50620 5850 50672 5856
rect 50160 5568 50212 5574
rect 50160 5510 50212 5516
rect 51080 5568 51132 5574
rect 51080 5510 51132 5516
rect 49332 4004 49384 4010
rect 49332 3946 49384 3952
rect 50172 3942 50200 5510
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 51092 5302 51120 5510
rect 51080 5296 51132 5302
rect 51080 5238 51132 5244
rect 52184 5024 52236 5030
rect 52184 4966 52236 4972
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 49620 3126 49648 3470
rect 49608 3120 49660 3126
rect 49608 3062 49660 3068
rect 50172 3058 50200 3878
rect 51170 3632 51226 3641
rect 51170 3567 51172 3576
rect 51224 3567 51226 3576
rect 51172 3538 51224 3544
rect 51538 3496 51594 3505
rect 51538 3431 51594 3440
rect 51552 3398 51580 3431
rect 51540 3392 51592 3398
rect 51540 3334 51592 3340
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 50160 3052 50212 3058
rect 50160 2994 50212 3000
rect 51552 2990 51580 3334
rect 52196 3058 52224 4966
rect 52184 3052 52236 3058
rect 52184 2994 52236 3000
rect 51540 2984 51592 2990
rect 51540 2926 51592 2932
rect 50160 2916 50212 2922
rect 50160 2858 50212 2864
rect 49056 2576 49108 2582
rect 49056 2518 49108 2524
rect 49424 2440 49476 2446
rect 49424 2382 49476 2388
rect 48872 2304 48924 2310
rect 48872 2246 48924 2252
rect 48884 1562 48912 2246
rect 48872 1556 48924 1562
rect 48872 1498 48924 1504
rect 49436 800 49464 2382
rect 49896 870 50016 898
rect 49896 800 49924 870
rect 46584 734 46796 762
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 49988 762 50016 870
rect 50172 762 50200 2858
rect 51356 2848 51408 2854
rect 51356 2790 51408 2796
rect 51264 2508 51316 2514
rect 51264 2450 51316 2456
rect 50896 2440 50948 2446
rect 51276 2417 51304 2450
rect 50896 2382 50948 2388
rect 51262 2408 51318 2417
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50908 800 50936 2382
rect 51262 2343 51318 2352
rect 51368 800 51396 2790
rect 52656 2514 52684 6598
rect 57152 3732 57204 3738
rect 57152 3674 57204 3680
rect 57164 3126 57192 3674
rect 58164 3528 58216 3534
rect 58164 3470 58216 3476
rect 57152 3120 57204 3126
rect 57152 3062 57204 3068
rect 55864 3052 55916 3058
rect 55864 2994 55916 3000
rect 55876 2961 55904 2994
rect 55862 2952 55918 2961
rect 55862 2887 55918 2896
rect 52828 2848 52880 2854
rect 52828 2790 52880 2796
rect 54300 2848 54352 2854
rect 54300 2790 54352 2796
rect 55772 2848 55824 2854
rect 55772 2790 55824 2796
rect 52644 2508 52696 2514
rect 52644 2450 52696 2456
rect 52368 2440 52420 2446
rect 52368 2382 52420 2388
rect 52380 800 52408 2382
rect 52840 800 52868 2790
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53012 2372 53064 2378
rect 53012 2314 53064 2320
rect 53024 1630 53052 2314
rect 53012 1624 53064 1630
rect 53012 1566 53064 1572
rect 53852 800 53880 2382
rect 54208 2372 54260 2378
rect 54208 2314 54260 2320
rect 54220 1766 54248 2314
rect 54208 1760 54260 1766
rect 54208 1702 54260 1708
rect 54312 800 54340 2790
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 55232 800 55260 2382
rect 55588 2372 55640 2378
rect 55588 2314 55640 2320
rect 55600 1834 55628 2314
rect 55588 1828 55640 1834
rect 55588 1770 55640 1776
rect 55784 800 55812 2790
rect 56692 2440 56744 2446
rect 56692 2382 56744 2388
rect 56704 800 56732 2382
rect 57060 2372 57112 2378
rect 57060 2314 57112 2320
rect 57072 1970 57100 2314
rect 57244 2304 57296 2310
rect 57244 2246 57296 2252
rect 57060 1964 57112 1970
rect 57060 1906 57112 1912
rect 57256 800 57284 2246
rect 58176 800 58204 3470
rect 59636 3188 59688 3194
rect 59636 3130 59688 3136
rect 58716 2848 58768 2854
rect 58716 2790 58768 2796
rect 58728 800 58756 2790
rect 59648 800 59676 3130
rect 49988 734 50200 762
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< via2 >>
rect 2962 41656 3018 41712
rect 2778 40024 2834 40080
rect 1582 39244 1584 39264
rect 1584 39244 1636 39264
rect 1636 39244 1638 39264
rect 1582 39208 1638 39244
rect 1582 38392 1638 38448
rect 1582 37612 1584 37632
rect 1584 37612 1636 37632
rect 1636 37612 1638 37632
rect 1582 37576 1638 37612
rect 1582 36644 1638 36680
rect 1582 36624 1584 36644
rect 1584 36624 1636 36644
rect 1636 36624 1638 36644
rect 1582 35808 1638 35864
rect 1582 34992 1638 35048
rect 1582 33804 1584 33824
rect 1584 33804 1636 33824
rect 1636 33804 1638 33824
rect 1582 33768 1638 33804
rect 1398 33360 1454 33416
rect 1582 32408 1638 32464
rect 1398 32000 1454 32056
rect 1582 31184 1638 31240
rect 3054 40840 3110 40896
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 1858 34584 1914 34640
rect 1398 29144 1454 29200
rect 1766 30776 1822 30832
rect 1582 29960 1638 30016
rect 1674 29588 1676 29608
rect 1676 29588 1728 29608
rect 1728 29588 1730 29608
rect 1674 29552 1730 29588
rect 1582 28736 1638 28792
rect 1582 27376 1638 27432
rect 1582 26188 1584 26208
rect 1584 26188 1636 26208
rect 1636 26188 1638 26208
rect 1582 26152 1638 26188
rect 1582 24928 1638 24984
rect 1490 24520 1546 24576
rect 1582 24112 1638 24168
rect 1858 28328 1914 28384
rect 1858 26968 1914 27024
rect 1858 25744 1914 25800
rect 1582 23704 1638 23760
rect 1398 23180 1454 23216
rect 1398 23160 1400 23180
rect 1400 23160 1452 23180
rect 1452 23160 1454 23180
rect 1582 22380 1584 22400
rect 1584 22380 1636 22400
rect 1636 22380 1638 22400
rect 1582 22344 1638 22380
rect 1858 21972 1860 21992
rect 1860 21972 1912 21992
rect 1912 21972 1914 21992
rect 1858 21936 1914 21972
rect 1582 21120 1638 21176
rect 1582 19896 1638 19952
rect 1398 17720 1454 17776
rect 1582 18536 1638 18592
rect 1858 19488 1914 19544
rect 1858 18128 1914 18184
rect 2318 34176 2374 34232
rect 2318 31592 2374 31648
rect 2318 30096 2374 30152
rect 2778 32952 2834 33008
rect 2594 30096 2650 30152
rect 3054 30368 3110 30424
rect 2870 25336 2926 25392
rect 1398 16088 1454 16144
rect 1582 15680 1638 15736
rect 1582 14864 1638 14920
rect 1398 14476 1454 14512
rect 1398 14456 1400 14476
rect 1400 14456 1452 14476
rect 1452 14456 1454 14476
rect 2226 19080 2282 19136
rect 2870 21528 2926 21584
rect 3054 20712 3110 20768
rect 2778 20304 2834 20360
rect 3974 27784 4030 27840
rect 3974 26560 4030 26616
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 3974 22752 4030 22808
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 2870 17312 2926 17368
rect 2686 17040 2742 17096
rect 3330 16904 3386 16960
rect 3974 16532 3976 16552
rect 3976 16532 4028 16552
rect 4028 16532 4030 16552
rect 3974 16496 4030 16532
rect 2318 13932 2374 13968
rect 2318 13912 2320 13932
rect 2320 13912 2372 13932
rect 2372 13912 2374 13932
rect 3974 15272 4030 15328
rect 1582 13504 1638 13560
rect 1858 13096 1914 13152
rect 1398 12688 1454 12744
rect 1582 12280 1638 12336
rect 1582 11464 1638 11520
rect 1582 11056 1638 11112
rect 1582 10240 1638 10296
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1766 8880 1822 8936
rect 1398 8064 1454 8120
rect 1582 7656 1638 7712
rect 2318 6840 2374 6896
rect 1398 6432 1454 6488
rect 1582 6060 1584 6080
rect 1584 6060 1636 6080
rect 1636 6060 1638 6080
rect 1582 6024 1638 6060
rect 3330 11872 3386 11928
rect 3054 10648 3110 10704
rect 2870 8472 2926 8528
rect 2962 7248 3018 7304
rect 1858 5616 1914 5672
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2962 4664 3018 4720
rect 2870 4256 2926 4312
rect 1858 3848 1914 3904
rect 1858 1808 1914 1864
rect 2686 3476 2688 3496
rect 2688 3476 2740 3496
rect 2740 3476 2742 3496
rect 2686 3440 2742 3476
rect 1306 584 1362 640
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3790 4120 3846 4176
rect 3146 1400 3202 1456
rect 3330 1028 3332 1048
rect 3332 1028 3384 1048
rect 3384 1028 3386 1048
rect 3330 992 3386 1028
rect 3698 2644 3754 2680
rect 3698 2624 3700 2644
rect 3700 2624 3752 2644
rect 3752 2624 3754 2644
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4066 3032 4122 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3882 2216 3938 2272
rect 5538 4140 5594 4176
rect 5538 4120 5540 4140
rect 5540 4120 5592 4140
rect 5592 4120 5594 4140
rect 6458 3440 6514 3496
rect 6918 3712 6974 3768
rect 2870 176 2926 232
rect 9310 17720 9366 17776
rect 9126 17620 9128 17640
rect 9128 17620 9180 17640
rect 9180 17620 9182 17640
rect 9126 17584 9182 17620
rect 9126 17040 9182 17096
rect 9494 17740 9550 17776
rect 9494 17720 9496 17740
rect 9496 17720 9548 17740
rect 9548 17720 9550 17740
rect 9494 17584 9550 17640
rect 10506 23432 10562 23488
rect 9770 14456 9826 14512
rect 9954 12824 10010 12880
rect 9678 12588 9680 12608
rect 9680 12588 9732 12608
rect 9732 12588 9734 12608
rect 9678 12552 9734 12588
rect 10230 12144 10286 12200
rect 9218 3596 9274 3632
rect 9218 3576 9220 3596
rect 9220 3576 9272 3596
rect 9272 3576 9274 3596
rect 9126 3440 9182 3496
rect 10506 12688 10562 12744
rect 10874 16652 10930 16688
rect 10874 16632 10876 16652
rect 10876 16632 10928 16652
rect 10928 16632 10930 16652
rect 10598 3476 10600 3496
rect 10600 3476 10652 3496
rect 10652 3476 10654 3496
rect 10598 3440 10654 3476
rect 12530 12552 12586 12608
rect 10874 3576 10930 3632
rect 12438 3712 12494 3768
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 14002 19080 14058 19136
rect 13818 16632 13874 16688
rect 13910 16224 13966 16280
rect 14646 16788 14702 16824
rect 14646 16768 14648 16788
rect 14648 16768 14700 16788
rect 14700 16768 14702 16788
rect 15290 15564 15346 15600
rect 15290 15544 15292 15564
rect 15292 15544 15344 15564
rect 15344 15544 15346 15564
rect 15198 2488 15254 2544
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19430 22072 19486 22128
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19430 21120 19486 21176
rect 17498 16108 17554 16144
rect 17498 16088 17500 16108
rect 17500 16088 17552 16108
rect 17552 16088 17554 16108
rect 19430 20848 19486 20904
rect 19614 20848 19670 20904
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19338 20304 19394 20360
rect 19522 20168 19578 20224
rect 19890 20340 19892 20360
rect 19892 20340 19944 20360
rect 19944 20340 19946 20360
rect 19890 20304 19946 20340
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19154 19080 19210 19136
rect 18510 16904 18566 16960
rect 18602 16768 18658 16824
rect 19706 18944 19762 19000
rect 20350 21956 20406 21992
rect 20350 21936 20352 21956
rect 20352 21936 20404 21956
rect 20404 21936 20406 21956
rect 20258 20168 20314 20224
rect 20626 22092 20682 22128
rect 20626 22072 20628 22092
rect 20628 22072 20680 22092
rect 20680 22072 20682 22092
rect 20626 20848 20682 20904
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20626 17484 20628 17504
rect 20628 17484 20680 17504
rect 20680 17484 20682 17504
rect 20626 17448 20682 17484
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 18878 16904 18934 16960
rect 18786 16224 18842 16280
rect 18694 16108 18750 16144
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 21730 17040 21786 17096
rect 18694 16088 18696 16108
rect 18696 16088 18748 16108
rect 18748 16088 18750 16108
rect 20258 15580 20260 15600
rect 20260 15580 20312 15600
rect 20312 15580 20314 15600
rect 20258 15544 20314 15580
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 21638 15036 21640 15056
rect 21640 15036 21692 15056
rect 21692 15036 21694 15056
rect 21638 15000 21694 15036
rect 21638 14900 21640 14920
rect 21640 14900 21692 14920
rect 21692 14900 21694 14920
rect 21638 14864 21694 14900
rect 20902 14728 20958 14784
rect 24122 20052 24178 20088
rect 24122 20032 24124 20052
rect 24124 20032 24176 20052
rect 24176 20032 24178 20052
rect 22282 17196 22338 17232
rect 22282 17176 22284 17196
rect 22284 17176 22336 17196
rect 22336 17176 22338 17196
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 18418 10648 18474 10704
rect 19982 13096 20038 13152
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19430 11192 19486 11248
rect 19338 10920 19394 10976
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19522 10684 19524 10704
rect 19524 10684 19576 10704
rect 19576 10684 19578 10704
rect 19522 10648 19578 10684
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19338 9424 19394 9480
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19890 6296 19946 6352
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20258 3884 20260 3904
rect 20260 3884 20312 3904
rect 20312 3884 20314 3904
rect 20258 3848 20314 3884
rect 19062 2488 19118 2544
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21638 13640 21694 13696
rect 22098 14728 22154 14784
rect 21638 11636 21640 11656
rect 21640 11636 21692 11656
rect 21692 11636 21694 11656
rect 21638 11600 21694 11636
rect 22282 15000 22338 15056
rect 22006 9460 22008 9480
rect 22008 9460 22060 9480
rect 22060 9460 22062 9480
rect 22006 9424 22062 9460
rect 22374 11600 22430 11656
rect 22650 11736 22706 11792
rect 21178 7792 21234 7848
rect 20994 6876 20996 6896
rect 20996 6876 21048 6896
rect 21048 6876 21050 6896
rect 20994 6840 21050 6876
rect 22282 6840 22338 6896
rect 25686 17448 25742 17504
rect 26054 17040 26110 17096
rect 24398 12552 24454 12608
rect 23478 9460 23480 9480
rect 23480 9460 23532 9480
rect 23532 9460 23534 9480
rect 23478 9424 23534 9460
rect 22006 3984 22062 4040
rect 23294 5072 23350 5128
rect 22190 4004 22246 4040
rect 22190 3984 22192 4004
rect 22192 3984 22244 4004
rect 22244 3984 22246 4004
rect 22098 3712 22154 3768
rect 22926 3576 22982 3632
rect 24582 5616 24638 5672
rect 24674 4120 24730 4176
rect 25410 3712 25466 3768
rect 28446 21936 28502 21992
rect 27526 17196 27582 17232
rect 27526 17176 27528 17196
rect 27528 17176 27580 17196
rect 27580 17176 27582 17196
rect 28906 20032 28962 20088
rect 28170 14864 28226 14920
rect 28170 13096 28226 13152
rect 26882 7828 26884 7848
rect 26884 7828 26936 7848
rect 26936 7828 26938 7848
rect 26882 7792 26938 7828
rect 26974 5636 27030 5672
rect 26974 5616 26976 5636
rect 26976 5616 27028 5636
rect 27028 5616 27030 5636
rect 26974 3848 27030 3904
rect 27802 6296 27858 6352
rect 27986 3576 28042 3632
rect 28814 19216 28870 19272
rect 28906 18944 28962 19000
rect 31114 21548 31170 21584
rect 31114 21528 31116 21548
rect 31116 21528 31168 21548
rect 31168 21528 31170 21548
rect 29182 19216 29238 19272
rect 28814 13640 28870 13696
rect 28538 11736 28594 11792
rect 29642 19216 29698 19272
rect 29550 18264 29606 18320
rect 28814 12552 28870 12608
rect 29734 6160 29790 6216
rect 30838 18400 30894 18456
rect 30286 13932 30342 13968
rect 30286 13912 30288 13932
rect 30288 13912 30340 13932
rect 30340 13912 30342 13932
rect 30010 6452 30066 6488
rect 30010 6432 30012 6452
rect 30012 6432 30064 6452
rect 30064 6432 30066 6452
rect 29826 3032 29882 3088
rect 32218 21528 32274 21584
rect 31390 14864 31446 14920
rect 31114 4564 31116 4584
rect 31116 4564 31168 4584
rect 31168 4564 31170 4584
rect 31114 4528 31170 4564
rect 31022 3188 31078 3224
rect 31022 3168 31024 3188
rect 31024 3168 31076 3188
rect 31076 3168 31078 3188
rect 31758 14900 31760 14920
rect 31760 14900 31812 14920
rect 31812 14900 31814 14920
rect 31758 14864 31814 14900
rect 32218 19252 32220 19272
rect 32220 19252 32272 19272
rect 32272 19252 32274 19272
rect 32218 19216 32274 19252
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 32862 21548 32918 21584
rect 32862 21528 32864 21548
rect 32864 21528 32916 21548
rect 32916 21528 32918 21548
rect 31758 9460 31760 9480
rect 31760 9460 31812 9480
rect 31812 9460 31814 9480
rect 31758 9424 31814 9460
rect 32402 9288 32458 9344
rect 32402 9036 32458 9072
rect 32402 9016 32404 9036
rect 32404 9016 32456 9036
rect 32456 9016 32458 9036
rect 31942 8880 31998 8936
rect 32034 8336 32090 8392
rect 31850 3032 31906 3088
rect 33138 16088 33194 16144
rect 33690 21548 33746 21584
rect 33690 21528 33692 21548
rect 33692 21528 33744 21548
rect 33744 21528 33746 21548
rect 33506 18284 33562 18320
rect 33506 18264 33508 18284
rect 33508 18264 33560 18284
rect 33560 18264 33562 18284
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 33690 13932 33746 13968
rect 33690 13912 33692 13932
rect 33692 13912 33744 13932
rect 33744 13912 33746 13932
rect 32862 8472 32918 8528
rect 33782 9460 33784 9480
rect 33784 9460 33836 9480
rect 33836 9460 33838 9480
rect 33782 9424 33838 9460
rect 33782 8744 33838 8800
rect 33322 4564 33324 4584
rect 33324 4564 33376 4584
rect 33376 4564 33378 4584
rect 33322 4528 33378 4564
rect 33598 5208 33654 5264
rect 34426 16124 34428 16144
rect 34428 16124 34480 16144
rect 34480 16124 34482 16144
rect 34426 16088 34482 16124
rect 34334 9052 34336 9072
rect 34336 9052 34388 9072
rect 34388 9052 34390 9072
rect 34334 9016 34390 9052
rect 34334 8744 34390 8800
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35806 21564 35808 21584
rect 35808 21564 35860 21584
rect 35860 21564 35862 21584
rect 35806 21528 35862 21564
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35530 9152 35586 9208
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34702 5788 34704 5808
rect 34704 5788 34756 5808
rect 34756 5788 34758 5808
rect 34702 5752 34758 5788
rect 35346 4936 35402 4992
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35254 4664 35310 4720
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35254 2932 35256 2952
rect 35256 2932 35308 2952
rect 35308 2932 35310 2952
rect 35254 2896 35310 2932
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 9424 35954 9480
rect 35806 8372 35808 8392
rect 35808 8372 35860 8392
rect 35860 8372 35862 8392
rect 35806 8336 35862 8372
rect 35806 5752 35862 5808
rect 35714 4664 35770 4720
rect 36634 18400 36690 18456
rect 36818 9424 36874 9480
rect 36082 5208 36138 5264
rect 36082 4936 36138 4992
rect 36726 3168 36782 3224
rect 37370 6432 37426 6488
rect 37830 8336 37886 8392
rect 37738 4528 37794 4584
rect 38198 8880 38254 8936
rect 39210 9444 39266 9480
rect 39210 9424 39212 9444
rect 39212 9424 39264 9444
rect 39264 9424 39266 9444
rect 38934 9152 38990 9208
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 40682 12180 40684 12200
rect 40684 12180 40736 12200
rect 40736 12180 40738 12200
rect 40682 12144 40738 12180
rect 41142 11736 41198 11792
rect 42522 11756 42578 11792
rect 42522 11736 42524 11756
rect 42524 11736 42576 11756
rect 42576 11736 42578 11756
rect 40038 8508 40040 8528
rect 40040 8508 40092 8528
rect 40092 8508 40094 8528
rect 40038 8472 40094 8508
rect 38290 6604 38292 6624
rect 38292 6604 38344 6624
rect 38344 6604 38346 6624
rect 38290 6568 38346 6604
rect 38566 6180 38622 6216
rect 38566 6160 38568 6180
rect 38568 6160 38620 6180
rect 38620 6160 38622 6180
rect 39394 6180 39450 6216
rect 39394 6160 39396 6180
rect 39396 6160 39448 6180
rect 39448 6160 39450 6180
rect 40958 8336 41014 8392
rect 38566 4140 38622 4176
rect 38566 4120 38568 4140
rect 38568 4120 38620 4140
rect 38620 4120 38622 4140
rect 41234 5752 41290 5808
rect 41694 6568 41750 6624
rect 44086 12144 44142 12200
rect 43350 5788 43352 5808
rect 43352 5788 43404 5808
rect 43404 5788 43406 5808
rect 43350 5752 43406 5788
rect 40866 4120 40922 4176
rect 39578 3168 39634 3224
rect 37922 2932 37924 2952
rect 37924 2932 37976 2952
rect 37976 2932 37978 2952
rect 37922 2896 37978 2932
rect 40866 3168 40922 3224
rect 41326 3712 41382 3768
rect 42154 3596 42210 3632
rect 42154 3576 42156 3596
rect 42156 3576 42208 3596
rect 42208 3576 42210 3596
rect 42798 3732 42854 3768
rect 42798 3712 42800 3732
rect 42800 3712 42852 3732
rect 42852 3712 42854 3732
rect 43442 3712 43498 3768
rect 42706 3168 42762 3224
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 45742 5072 45798 5128
rect 45834 4140 45890 4176
rect 45834 4120 45836 4140
rect 45836 4120 45888 4140
rect 45888 4120 45890 4140
rect 45926 3476 45928 3496
rect 45928 3476 45980 3496
rect 45980 3476 45982 3496
rect 45926 3440 45982 3476
rect 47490 6160 47546 6216
rect 46846 4140 46902 4176
rect 46846 4120 46848 4140
rect 46848 4120 46900 4140
rect 46900 4120 46902 4140
rect 47582 3732 47638 3768
rect 47582 3712 47584 3732
rect 47584 3712 47636 3732
rect 47636 3712 47638 3732
rect 47582 3596 47638 3632
rect 47582 3576 47584 3596
rect 47584 3576 47636 3596
rect 47636 3576 47638 3596
rect 47214 3460 47270 3496
rect 47214 3440 47216 3460
rect 47216 3440 47268 3460
rect 47268 3440 47270 3460
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 47858 3476 47860 3496
rect 47860 3476 47912 3496
rect 47912 3476 47914 3496
rect 47858 3440 47914 3476
rect 48502 3596 48558 3632
rect 48502 3576 48504 3596
rect 48504 3576 48556 3596
rect 48556 3576 48558 3596
rect 48870 3476 48872 3496
rect 48872 3476 48924 3496
rect 48924 3476 48926 3496
rect 48870 3440 48926 3476
rect 48778 2896 48834 2952
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 51170 3596 51226 3632
rect 51170 3576 51172 3596
rect 51172 3576 51224 3596
rect 51224 3576 51226 3596
rect 51538 3440 51594 3496
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 51262 2352 51318 2408
rect 55862 2896 55918 2952
<< metal3 >>
rect 0 41714 800 41744
rect 2957 41714 3023 41717
rect 0 41712 3023 41714
rect 0 41656 2962 41712
rect 3018 41656 3023 41712
rect 0 41654 3023 41656
rect 0 41624 800 41654
rect 2957 41651 3023 41654
rect 0 41216 800 41336
rect 0 40898 800 40928
rect 3049 40898 3115 40901
rect 0 40896 3115 40898
rect 0 40840 3054 40896
rect 3110 40840 3115 40896
rect 0 40838 3115 40840
rect 0 40808 800 40838
rect 3049 40835 3115 40838
rect 0 40400 800 40520
rect 0 40082 800 40112
rect 2773 40082 2839 40085
rect 0 40080 2839 40082
rect 0 40024 2778 40080
rect 2834 40024 2839 40080
rect 0 40022 2839 40024
rect 0 39992 800 40022
rect 2773 40019 2839 40022
rect 4208 39744 4528 39745
rect 0 39584 800 39704
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39266 800 39296
rect 1577 39266 1643 39269
rect 0 39264 1643 39266
rect 0 39208 1582 39264
rect 1638 39208 1643 39264
rect 0 39206 1643 39208
rect 0 39176 800 39206
rect 1577 39203 1643 39206
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 50288 39200 50608 39201
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 39135 50608 39136
rect 0 38768 800 38888
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38450 800 38480
rect 1577 38450 1643 38453
rect 0 38448 1643 38450
rect 0 38392 1582 38448
rect 1638 38392 1643 38448
rect 0 38390 1643 38392
rect 0 38360 800 38390
rect 1577 38387 1643 38390
rect 19568 38112 19888 38113
rect 0 37952 800 38072
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 50288 38112 50608 38113
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 38047 50608 38048
rect 0 37634 800 37664
rect 1577 37634 1643 37637
rect 0 37632 1643 37634
rect 0 37576 1582 37632
rect 1638 37576 1643 37632
rect 0 37574 1643 37576
rect 0 37544 800 37574
rect 1577 37571 1643 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 0 37000 800 37120
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36184 800 36304
rect 19568 35936 19888 35937
rect 0 35866 800 35896
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 0 35368 800 35488
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 0 34642 800 34672
rect 1853 34642 1919 34645
rect 0 34640 1919 34642
rect 0 34584 1858 34640
rect 1914 34584 1919 34640
rect 0 34582 1919 34584
rect 0 34552 800 34582
rect 1853 34579 1919 34582
rect 4208 34304 4528 34305
rect 0 34234 800 34264
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 2313 34234 2379 34237
rect 0 34232 2379 34234
rect 0 34176 2318 34232
rect 2374 34176 2379 34232
rect 0 34174 2379 34176
rect 0 34144 800 34174
rect 2313 34171 2379 34174
rect 0 33826 800 33856
rect 1577 33826 1643 33829
rect 0 33824 1643 33826
rect 0 33768 1582 33824
rect 1638 33768 1643 33824
rect 0 33766 1643 33768
rect 0 33736 800 33766
rect 1577 33763 1643 33766
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 0 33418 800 33448
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33328 800 33358
rect 1393 33355 1459 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 33010 800 33040
rect 2773 33010 2839 33013
rect 0 33008 2839 33010
rect 0 32952 2778 33008
rect 2834 32952 2839 33008
rect 0 32950 2839 32952
rect 0 32920 800 32950
rect 2773 32947 2839 32950
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 1393 32058 1459 32061
rect 0 32056 1459 32058
rect 0 32000 1398 32056
rect 1454 32000 1459 32056
rect 0 31998 1459 32000
rect 0 31968 800 31998
rect 1393 31995 1459 31998
rect 0 31650 800 31680
rect 2313 31650 2379 31653
rect 0 31648 2379 31650
rect 0 31592 2318 31648
rect 2374 31592 2379 31648
rect 0 31590 2379 31592
rect 0 31560 800 31590
rect 2313 31587 2379 31590
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31242 800 31272
rect 1577 31242 1643 31245
rect 0 31240 1643 31242
rect 0 31184 1582 31240
rect 1638 31184 1643 31240
rect 0 31182 1643 31184
rect 0 31152 800 31182
rect 1577 31179 1643 31182
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 0 30834 800 30864
rect 1761 30834 1827 30837
rect 0 30832 1827 30834
rect 0 30776 1766 30832
rect 1822 30776 1827 30832
rect 0 30774 1827 30776
rect 0 30744 800 30774
rect 1761 30771 1827 30774
rect 19568 30496 19888 30497
rect 0 30426 800 30456
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 3049 30426 3115 30429
rect 0 30424 3115 30426
rect 0 30368 3054 30424
rect 3110 30368 3115 30424
rect 0 30366 3115 30368
rect 0 30336 800 30366
rect 3049 30363 3115 30366
rect 2313 30154 2379 30157
rect 2589 30154 2655 30157
rect 2313 30152 2655 30154
rect 2313 30096 2318 30152
rect 2374 30096 2594 30152
rect 2650 30096 2655 30152
rect 2313 30094 2655 30096
rect 2313 30091 2379 30094
rect 2589 30091 2655 30094
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 0 29610 800 29640
rect 1669 29610 1735 29613
rect 0 29608 1735 29610
rect 0 29552 1674 29608
rect 1730 29552 1735 29608
rect 0 29550 1735 29552
rect 0 29520 800 29550
rect 1669 29547 1735 29550
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 0 29202 800 29232
rect 1393 29202 1459 29205
rect 0 29200 1459 29202
rect 0 29144 1398 29200
rect 1454 29144 1459 29200
rect 0 29142 1459 29144
rect 0 29112 800 29142
rect 1393 29139 1459 29142
rect 4208 28864 4528 28865
rect 0 28794 800 28824
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 1577 28794 1643 28797
rect 0 28792 1643 28794
rect 0 28736 1582 28792
rect 1638 28736 1643 28792
rect 0 28734 1643 28736
rect 0 28704 800 28734
rect 1577 28731 1643 28734
rect 0 28386 800 28416
rect 1853 28386 1919 28389
rect 0 28384 1919 28386
rect 0 28328 1858 28384
rect 1914 28328 1919 28384
rect 0 28326 1919 28328
rect 0 28296 800 28326
rect 1853 28323 1919 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 0 27842 800 27872
rect 3969 27842 4035 27845
rect 0 27840 4035 27842
rect 0 27784 3974 27840
rect 4030 27784 4035 27840
rect 0 27782 4035 27784
rect 0 27752 800 27782
rect 3969 27779 4035 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 0 27026 800 27056
rect 1853 27026 1919 27029
rect 0 27024 1919 27026
rect 0 26968 1858 27024
rect 1914 26968 1919 27024
rect 0 26966 1919 26968
rect 0 26936 800 26966
rect 1853 26963 1919 26966
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 3969 26618 4035 26621
rect 0 26616 4035 26618
rect 0 26560 3974 26616
rect 4030 26560 4035 26616
rect 0 26558 4035 26560
rect 0 26528 800 26558
rect 3969 26555 4035 26558
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 0 25802 800 25832
rect 1853 25802 1919 25805
rect 0 25800 1919 25802
rect 0 25744 1858 25800
rect 1914 25744 1919 25800
rect 0 25742 1919 25744
rect 0 25712 800 25742
rect 1853 25739 1919 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25394 800 25424
rect 2865 25394 2931 25397
rect 0 25392 2931 25394
rect 0 25336 2870 25392
rect 2926 25336 2931 25392
rect 0 25334 2931 25336
rect 0 25304 800 25334
rect 2865 25331 2931 25334
rect 19568 25056 19888 25057
rect 0 24986 800 25016
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 0 24578 800 24608
rect 1485 24578 1551 24581
rect 0 24576 1551 24578
rect 0 24520 1490 24576
rect 1546 24520 1551 24576
rect 0 24518 1551 24520
rect 0 24488 800 24518
rect 1485 24515 1551 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 0 23762 800 23792
rect 1577 23762 1643 23765
rect 0 23760 1643 23762
rect 0 23704 1582 23760
rect 1638 23704 1643 23760
rect 0 23702 1643 23704
rect 0 23672 800 23702
rect 1577 23699 1643 23702
rect 10501 23492 10567 23493
rect 10501 23488 10548 23492
rect 10612 23490 10618 23492
rect 10501 23432 10506 23488
rect 10501 23428 10548 23432
rect 10612 23430 10658 23490
rect 10612 23428 10618 23430
rect 10501 23427 10567 23428
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 19568 22880 19888 22881
rect 0 22810 800 22840
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 3969 22810 4035 22813
rect 0 22808 4035 22810
rect 0 22752 3974 22808
rect 4030 22752 4035 22808
rect 0 22750 4035 22752
rect 0 22720 800 22750
rect 3969 22747 4035 22750
rect 0 22402 800 22432
rect 1577 22402 1643 22405
rect 0 22400 1643 22402
rect 0 22344 1582 22400
rect 1638 22344 1643 22400
rect 0 22342 1643 22344
rect 0 22312 800 22342
rect 1577 22339 1643 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 19425 22130 19491 22133
rect 20621 22130 20687 22133
rect 19425 22128 20687 22130
rect 19425 22072 19430 22128
rect 19486 22072 20626 22128
rect 20682 22072 20687 22128
rect 19425 22070 20687 22072
rect 19425 22067 19491 22070
rect 20621 22067 20687 22070
rect 0 21994 800 22024
rect 1853 21994 1919 21997
rect 0 21992 1919 21994
rect 0 21936 1858 21992
rect 1914 21936 1919 21992
rect 0 21934 1919 21936
rect 0 21904 800 21934
rect 1853 21931 1919 21934
rect 20345 21994 20411 21997
rect 28441 21994 28507 21997
rect 20345 21992 28507 21994
rect 20345 21936 20350 21992
rect 20406 21936 28446 21992
rect 28502 21936 28507 21992
rect 20345 21934 28507 21936
rect 20345 21931 20411 21934
rect 28441 21931 28507 21934
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 0 21586 800 21616
rect 2865 21586 2931 21589
rect 0 21584 2931 21586
rect 0 21528 2870 21584
rect 2926 21528 2931 21584
rect 0 21526 2931 21528
rect 0 21496 800 21526
rect 2865 21523 2931 21526
rect 31109 21586 31175 21589
rect 32213 21586 32279 21589
rect 32857 21586 32923 21589
rect 31109 21584 32923 21586
rect 31109 21528 31114 21584
rect 31170 21528 32218 21584
rect 32274 21528 32862 21584
rect 32918 21528 32923 21584
rect 31109 21526 32923 21528
rect 31109 21523 31175 21526
rect 32213 21523 32279 21526
rect 32857 21523 32923 21526
rect 33685 21586 33751 21589
rect 35801 21586 35867 21589
rect 33685 21584 35867 21586
rect 33685 21528 33690 21584
rect 33746 21528 35806 21584
rect 35862 21528 35867 21584
rect 33685 21526 35867 21528
rect 33685 21523 33751 21526
rect 35801 21523 35867 21526
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 1577 21178 1643 21181
rect 19425 21178 19491 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 19382 21176 19491 21178
rect 19382 21120 19430 21176
rect 19486 21120 19491 21176
rect 19382 21115 19491 21120
rect 19382 20909 19442 21115
rect 19382 20904 19491 20909
rect 19382 20848 19430 20904
rect 19486 20848 19491 20904
rect 19382 20846 19491 20848
rect 19425 20843 19491 20846
rect 19609 20906 19675 20909
rect 20621 20906 20687 20909
rect 19609 20904 20687 20906
rect 19609 20848 19614 20904
rect 19670 20848 20626 20904
rect 20682 20848 20687 20904
rect 19609 20846 20687 20848
rect 19609 20843 19675 20846
rect 20621 20843 20687 20846
rect 0 20770 800 20800
rect 3049 20770 3115 20773
rect 0 20768 3115 20770
rect 0 20712 3054 20768
rect 3110 20712 3115 20768
rect 0 20710 3115 20712
rect 0 20680 800 20710
rect 3049 20707 3115 20710
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 19333 20362 19399 20365
rect 19885 20362 19951 20365
rect 19333 20360 19951 20362
rect 19333 20304 19338 20360
rect 19394 20304 19890 20360
rect 19946 20304 19951 20360
rect 19333 20302 19951 20304
rect 19333 20299 19399 20302
rect 19885 20299 19951 20302
rect 19517 20226 19583 20229
rect 20253 20226 20319 20229
rect 19517 20224 20319 20226
rect 19517 20168 19522 20224
rect 19578 20168 20258 20224
rect 20314 20168 20319 20224
rect 19517 20166 20319 20168
rect 19517 20163 19583 20166
rect 20253 20163 20319 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 24117 20090 24183 20093
rect 28901 20090 28967 20093
rect 24117 20088 28967 20090
rect 24117 20032 24122 20088
rect 24178 20032 28906 20088
rect 28962 20032 28967 20088
rect 24117 20030 28967 20032
rect 24117 20027 24183 20030
rect 28901 20027 28967 20030
rect 0 19954 800 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 800 19894
rect 1577 19891 1643 19894
rect 19568 19616 19888 19617
rect 0 19546 800 19576
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 1853 19546 1919 19549
rect 0 19544 1919 19546
rect 0 19488 1858 19544
rect 1914 19488 1919 19544
rect 0 19486 1919 19488
rect 0 19456 800 19486
rect 1853 19483 1919 19486
rect 28809 19274 28875 19277
rect 29177 19274 29243 19277
rect 29637 19274 29703 19277
rect 32213 19274 32279 19277
rect 28809 19272 32279 19274
rect 28809 19216 28814 19272
rect 28870 19216 29182 19272
rect 29238 19216 29642 19272
rect 29698 19216 32218 19272
rect 32274 19216 32279 19272
rect 28809 19214 32279 19216
rect 28809 19211 28875 19214
rect 29177 19211 29243 19214
rect 29637 19211 29703 19214
rect 32213 19211 32279 19214
rect 0 19138 800 19168
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 19048 800 19078
rect 2221 19075 2287 19078
rect 13997 19138 14063 19141
rect 19149 19138 19215 19141
rect 13997 19136 19215 19138
rect 13997 19080 14002 19136
rect 14058 19080 19154 19136
rect 19210 19080 19215 19136
rect 13997 19078 19215 19080
rect 13997 19075 14063 19078
rect 19149 19075 19215 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19701 19002 19767 19005
rect 28901 19002 28967 19005
rect 19701 19000 28967 19002
rect 19701 18944 19706 19000
rect 19762 18944 28906 19000
rect 28962 18944 28967 19000
rect 19701 18942 28967 18944
rect 19701 18939 19767 18942
rect 28901 18939 28967 18942
rect 0 18594 800 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 800 18534
rect 1577 18531 1643 18534
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 30833 18458 30899 18461
rect 36629 18458 36695 18461
rect 30833 18456 36695 18458
rect 30833 18400 30838 18456
rect 30894 18400 36634 18456
rect 36690 18400 36695 18456
rect 30833 18398 36695 18400
rect 30833 18395 30899 18398
rect 36629 18395 36695 18398
rect 29545 18322 29611 18325
rect 33501 18322 33567 18325
rect 29545 18320 33567 18322
rect 29545 18264 29550 18320
rect 29606 18264 33506 18320
rect 33562 18264 33567 18320
rect 29545 18262 33567 18264
rect 29545 18259 29611 18262
rect 33501 18259 33567 18262
rect 0 18186 800 18216
rect 1853 18186 1919 18189
rect 0 18184 1919 18186
rect 0 18128 1858 18184
rect 1914 18128 1919 18184
rect 0 18126 1919 18128
rect 0 18096 800 18126
rect 1853 18123 1919 18126
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 9305 17778 9371 17781
rect 9489 17778 9555 17781
rect 9305 17776 9555 17778
rect 9305 17720 9310 17776
rect 9366 17720 9494 17776
rect 9550 17720 9555 17776
rect 9305 17718 9555 17720
rect 9305 17715 9371 17718
rect 9489 17715 9555 17718
rect 9121 17642 9187 17645
rect 9489 17642 9555 17645
rect 9121 17640 9555 17642
rect 9121 17584 9126 17640
rect 9182 17584 9494 17640
rect 9550 17584 9555 17640
rect 9121 17582 9555 17584
rect 9121 17579 9187 17582
rect 9489 17579 9555 17582
rect 20621 17506 20687 17509
rect 25681 17506 25747 17509
rect 20621 17504 25747 17506
rect 20621 17448 20626 17504
rect 20682 17448 25686 17504
rect 25742 17448 25747 17504
rect 20621 17446 25747 17448
rect 20621 17443 20687 17446
rect 25681 17443 25747 17446
rect 19568 17440 19888 17441
rect 0 17370 800 17400
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 2865 17370 2931 17373
rect 0 17368 2931 17370
rect 0 17312 2870 17368
rect 2926 17312 2931 17368
rect 0 17310 2931 17312
rect 0 17280 800 17310
rect 2865 17307 2931 17310
rect 22277 17234 22343 17237
rect 27521 17234 27587 17237
rect 22277 17232 27587 17234
rect 22277 17176 22282 17232
rect 22338 17176 27526 17232
rect 27582 17176 27587 17232
rect 22277 17174 27587 17176
rect 22277 17171 22343 17174
rect 27521 17171 27587 17174
rect 2681 17098 2747 17101
rect 9121 17098 9187 17101
rect 2681 17096 9187 17098
rect 2681 17040 2686 17096
rect 2742 17040 9126 17096
rect 9182 17040 9187 17096
rect 2681 17038 9187 17040
rect 2681 17035 2747 17038
rect 9121 17035 9187 17038
rect 21725 17098 21791 17101
rect 26049 17098 26115 17101
rect 21725 17096 26115 17098
rect 21725 17040 21730 17096
rect 21786 17040 26054 17096
rect 26110 17040 26115 17096
rect 21725 17038 26115 17040
rect 21725 17035 21791 17038
rect 26049 17035 26115 17038
rect 0 16962 800 16992
rect 3325 16962 3391 16965
rect 0 16960 3391 16962
rect 0 16904 3330 16960
rect 3386 16904 3391 16960
rect 0 16902 3391 16904
rect 0 16872 800 16902
rect 3325 16899 3391 16902
rect 18505 16962 18571 16965
rect 18873 16962 18939 16965
rect 18505 16960 18939 16962
rect 18505 16904 18510 16960
rect 18566 16904 18878 16960
rect 18934 16904 18939 16960
rect 18505 16902 18939 16904
rect 18505 16899 18571 16902
rect 18873 16899 18939 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 14641 16826 14707 16829
rect 18597 16826 18663 16829
rect 14641 16824 18663 16826
rect 14641 16768 14646 16824
rect 14702 16768 18602 16824
rect 18658 16768 18663 16824
rect 14641 16766 18663 16768
rect 14641 16763 14707 16766
rect 18597 16763 18663 16766
rect 10869 16690 10935 16693
rect 13813 16690 13879 16693
rect 10869 16688 13879 16690
rect 10869 16632 10874 16688
rect 10930 16632 13818 16688
rect 13874 16632 13879 16688
rect 10869 16630 13879 16632
rect 10869 16627 10935 16630
rect 13813 16627 13879 16630
rect 0 16554 800 16584
rect 3969 16554 4035 16557
rect 0 16552 4035 16554
rect 0 16496 3974 16552
rect 4030 16496 4035 16552
rect 0 16494 4035 16496
rect 0 16464 800 16494
rect 3969 16491 4035 16494
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 13905 16282 13971 16285
rect 18781 16282 18847 16285
rect 13905 16280 18847 16282
rect 13905 16224 13910 16280
rect 13966 16224 18786 16280
rect 18842 16224 18847 16280
rect 13905 16222 18847 16224
rect 13905 16219 13971 16222
rect 18781 16219 18847 16222
rect 0 16146 800 16176
rect 1393 16146 1459 16149
rect 0 16144 1459 16146
rect 0 16088 1398 16144
rect 1454 16088 1459 16144
rect 0 16086 1459 16088
rect 0 16056 800 16086
rect 1393 16083 1459 16086
rect 17493 16146 17559 16149
rect 18689 16146 18755 16149
rect 17493 16144 18755 16146
rect 17493 16088 17498 16144
rect 17554 16088 18694 16144
rect 18750 16088 18755 16144
rect 17493 16086 18755 16088
rect 17493 16083 17559 16086
rect 18689 16083 18755 16086
rect 33133 16146 33199 16149
rect 34421 16146 34487 16149
rect 33133 16144 34487 16146
rect 33133 16088 33138 16144
rect 33194 16088 34426 16144
rect 34482 16088 34487 16144
rect 33133 16086 34487 16088
rect 33133 16083 33199 16086
rect 34421 16083 34487 16086
rect 4208 15808 4528 15809
rect 0 15738 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 1577 15738 1643 15741
rect 0 15736 1643 15738
rect 0 15680 1582 15736
rect 1638 15680 1643 15736
rect 0 15678 1643 15680
rect 0 15648 800 15678
rect 1577 15675 1643 15678
rect 15285 15602 15351 15605
rect 20253 15602 20319 15605
rect 15285 15600 20319 15602
rect 15285 15544 15290 15600
rect 15346 15544 20258 15600
rect 20314 15544 20319 15600
rect 15285 15542 20319 15544
rect 15285 15539 15351 15542
rect 20253 15539 20319 15542
rect 0 15330 800 15360
rect 3969 15330 4035 15333
rect 0 15328 4035 15330
rect 0 15272 3974 15328
rect 4030 15272 4035 15328
rect 0 15270 4035 15272
rect 0 15240 800 15270
rect 3969 15267 4035 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 21633 15058 21699 15061
rect 22277 15058 22343 15061
rect 21633 15056 22343 15058
rect 21633 15000 21638 15056
rect 21694 15000 22282 15056
rect 22338 15000 22343 15056
rect 21633 14998 22343 15000
rect 21633 14995 21699 14998
rect 22277 14995 22343 14998
rect 0 14922 800 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 800 14862
rect 1577 14859 1643 14862
rect 21633 14922 21699 14925
rect 28165 14922 28231 14925
rect 21633 14920 28231 14922
rect 21633 14864 21638 14920
rect 21694 14864 28170 14920
rect 28226 14864 28231 14920
rect 21633 14862 28231 14864
rect 21633 14859 21699 14862
rect 28165 14859 28231 14862
rect 31385 14922 31451 14925
rect 31753 14922 31819 14925
rect 31385 14920 31819 14922
rect 31385 14864 31390 14920
rect 31446 14864 31758 14920
rect 31814 14864 31819 14920
rect 31385 14862 31819 14864
rect 31385 14859 31451 14862
rect 31753 14859 31819 14862
rect 20897 14786 20963 14789
rect 22093 14786 22159 14789
rect 20897 14784 22159 14786
rect 20897 14728 20902 14784
rect 20958 14728 22098 14784
rect 22154 14728 22159 14784
rect 20897 14726 22159 14728
rect 20897 14723 20963 14726
rect 22093 14723 22159 14726
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14514 800 14544
rect 1393 14514 1459 14517
rect 9765 14516 9831 14517
rect 9765 14514 9812 14516
rect 0 14512 1459 14514
rect 0 14456 1398 14512
rect 1454 14456 1459 14512
rect 0 14454 1459 14456
rect 9720 14512 9812 14514
rect 9720 14456 9770 14512
rect 9720 14454 9812 14456
rect 0 14424 800 14454
rect 1393 14451 1459 14454
rect 9765 14452 9812 14454
rect 9876 14452 9882 14516
rect 9765 14451 9831 14452
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 0 13970 800 14000
rect 2313 13970 2379 13973
rect 0 13968 2379 13970
rect 0 13912 2318 13968
rect 2374 13912 2379 13968
rect 0 13910 2379 13912
rect 0 13880 800 13910
rect 2313 13907 2379 13910
rect 30281 13970 30347 13973
rect 33685 13970 33751 13973
rect 30281 13968 33751 13970
rect 30281 13912 30286 13968
rect 30342 13912 33690 13968
rect 33746 13912 33751 13968
rect 30281 13910 33751 13912
rect 30281 13907 30347 13910
rect 33685 13907 33751 13910
rect 21633 13698 21699 13701
rect 28809 13698 28875 13701
rect 21633 13696 28875 13698
rect 21633 13640 21638 13696
rect 21694 13640 28814 13696
rect 28870 13640 28875 13696
rect 21633 13638 28875 13640
rect 21633 13635 21699 13638
rect 28809 13635 28875 13638
rect 4208 13632 4528 13633
rect 0 13562 800 13592
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 0 13154 800 13184
rect 1853 13154 1919 13157
rect 0 13152 1919 13154
rect 0 13096 1858 13152
rect 1914 13096 1919 13152
rect 0 13094 1919 13096
rect 0 13064 800 13094
rect 1853 13091 1919 13094
rect 19977 13154 20043 13157
rect 28165 13154 28231 13157
rect 19977 13152 28231 13154
rect 19977 13096 19982 13152
rect 20038 13096 28170 13152
rect 28226 13096 28231 13152
rect 19977 13094 28231 13096
rect 19977 13091 20043 13094
rect 28165 13091 28231 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 9949 12882 10015 12885
rect 9949 12880 10058 12882
rect 9949 12824 9954 12880
rect 10010 12824 10058 12880
rect 9949 12819 10058 12824
rect 0 12746 800 12776
rect 1393 12746 1459 12749
rect 0 12744 1459 12746
rect 0 12688 1398 12744
rect 1454 12688 1459 12744
rect 0 12686 1459 12688
rect 9998 12746 10058 12819
rect 10501 12746 10567 12749
rect 9998 12744 10567 12746
rect 9998 12688 10506 12744
rect 10562 12688 10567 12744
rect 9998 12686 10567 12688
rect 0 12656 800 12686
rect 1393 12683 1459 12686
rect 10501 12683 10567 12686
rect 9673 12610 9739 12613
rect 12525 12610 12591 12613
rect 9673 12608 12591 12610
rect 9673 12552 9678 12608
rect 9734 12552 12530 12608
rect 12586 12552 12591 12608
rect 9673 12550 12591 12552
rect 9673 12547 9739 12550
rect 12525 12547 12591 12550
rect 24393 12610 24459 12613
rect 28809 12610 28875 12613
rect 24393 12608 28875 12610
rect 24393 12552 24398 12608
rect 24454 12552 28814 12608
rect 28870 12552 28875 12608
rect 24393 12550 28875 12552
rect 24393 12547 24459 12550
rect 28809 12547 28875 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 9806 12140 9812 12204
rect 9876 12202 9882 12204
rect 10225 12202 10291 12205
rect 9876 12200 10291 12202
rect 9876 12144 10230 12200
rect 10286 12144 10291 12200
rect 9876 12142 10291 12144
rect 9876 12140 9882 12142
rect 10225 12139 10291 12142
rect 40677 12202 40743 12205
rect 44081 12202 44147 12205
rect 40677 12200 44147 12202
rect 40677 12144 40682 12200
rect 40738 12144 44086 12200
rect 44142 12144 44147 12200
rect 40677 12142 44147 12144
rect 40677 12139 40743 12142
rect 44081 12139 44147 12142
rect 19568 12000 19888 12001
rect 0 11930 800 11960
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 3325 11930 3391 11933
rect 0 11928 3391 11930
rect 0 11872 3330 11928
rect 3386 11872 3391 11928
rect 0 11870 3391 11872
rect 0 11840 800 11870
rect 3325 11867 3391 11870
rect 22645 11794 22711 11797
rect 28533 11794 28599 11797
rect 22645 11792 28599 11794
rect 22645 11736 22650 11792
rect 22706 11736 28538 11792
rect 28594 11736 28599 11792
rect 22645 11734 28599 11736
rect 22645 11731 22711 11734
rect 28533 11731 28599 11734
rect 41137 11794 41203 11797
rect 42517 11794 42583 11797
rect 41137 11792 42583 11794
rect 41137 11736 41142 11792
rect 41198 11736 42522 11792
rect 42578 11736 42583 11792
rect 41137 11734 42583 11736
rect 41137 11731 41203 11734
rect 42517 11731 42583 11734
rect 21633 11658 21699 11661
rect 22369 11658 22435 11661
rect 21633 11656 22435 11658
rect 21633 11600 21638 11656
rect 21694 11600 22374 11656
rect 22430 11600 22435 11656
rect 21633 11598 22435 11600
rect 21633 11595 21699 11598
rect 22369 11595 22435 11598
rect 0 11522 800 11552
rect 1577 11522 1643 11525
rect 0 11520 1643 11522
rect 0 11464 1582 11520
rect 1638 11464 1643 11520
rect 0 11462 1643 11464
rect 0 11432 800 11462
rect 1577 11459 1643 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 19425 11250 19491 11253
rect 19382 11248 19491 11250
rect 19382 11192 19430 11248
rect 19486 11192 19491 11248
rect 19382 11187 19491 11192
rect 0 11114 800 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 800 11054
rect 1577 11051 1643 11054
rect 19382 10981 19442 11187
rect 19333 10976 19442 10981
rect 19333 10920 19338 10976
rect 19394 10920 19442 10976
rect 19333 10918 19442 10920
rect 19333 10915 19399 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 0 10706 800 10736
rect 3049 10706 3115 10709
rect 0 10704 3115 10706
rect 0 10648 3054 10704
rect 3110 10648 3115 10704
rect 0 10646 3115 10648
rect 0 10616 800 10646
rect 3049 10643 3115 10646
rect 18413 10706 18479 10709
rect 19517 10706 19583 10709
rect 18413 10704 19583 10706
rect 18413 10648 18418 10704
rect 18474 10648 19522 10704
rect 19578 10648 19583 10704
rect 18413 10646 19583 10648
rect 18413 10643 18479 10646
rect 19517 10643 19583 10646
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 0 9800 800 9920
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 19333 9482 19399 9485
rect 22001 9482 22067 9485
rect 23473 9482 23539 9485
rect 19333 9480 23539 9482
rect 19333 9424 19338 9480
rect 19394 9424 22006 9480
rect 22062 9424 23478 9480
rect 23534 9424 23539 9480
rect 19333 9422 23539 9424
rect 19333 9419 19399 9422
rect 22001 9419 22067 9422
rect 23473 9419 23539 9422
rect 31753 9482 31819 9485
rect 33777 9482 33843 9485
rect 35893 9482 35959 9485
rect 31753 9480 33843 9482
rect 31753 9424 31758 9480
rect 31814 9424 33782 9480
rect 33838 9424 33843 9480
rect 31753 9422 33843 9424
rect 31753 9419 31819 9422
rect 33777 9419 33843 9422
rect 33918 9480 35959 9482
rect 33918 9424 35898 9480
rect 35954 9424 35959 9480
rect 33918 9422 35959 9424
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 32397 9346 32463 9349
rect 33918 9346 33978 9422
rect 35893 9419 35959 9422
rect 36813 9482 36879 9485
rect 39205 9482 39271 9485
rect 36813 9480 39271 9482
rect 36813 9424 36818 9480
rect 36874 9424 39210 9480
rect 39266 9424 39271 9480
rect 36813 9422 39271 9424
rect 36813 9419 36879 9422
rect 39205 9419 39271 9422
rect 32397 9344 33978 9346
rect 32397 9288 32402 9344
rect 32458 9288 33978 9344
rect 32397 9286 33978 9288
rect 32397 9283 32463 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 35525 9210 35591 9213
rect 38929 9210 38995 9213
rect 35525 9208 38995 9210
rect 35525 9152 35530 9208
rect 35586 9152 38934 9208
rect 38990 9152 38995 9208
rect 35525 9150 38995 9152
rect 35525 9147 35591 9150
rect 38929 9147 38995 9150
rect 32397 9074 32463 9077
rect 34329 9074 34395 9077
rect 32397 9072 34395 9074
rect 32397 9016 32402 9072
rect 32458 9016 34334 9072
rect 34390 9016 34395 9072
rect 32397 9014 34395 9016
rect 32397 9011 32463 9014
rect 34329 9011 34395 9014
rect 0 8938 800 8968
rect 1761 8938 1827 8941
rect 0 8936 1827 8938
rect 0 8880 1766 8936
rect 1822 8880 1827 8936
rect 0 8878 1827 8880
rect 0 8848 800 8878
rect 1761 8875 1827 8878
rect 31937 8938 32003 8941
rect 38193 8938 38259 8941
rect 31937 8936 38259 8938
rect 31937 8880 31942 8936
rect 31998 8880 38198 8936
rect 38254 8880 38259 8936
rect 31937 8878 38259 8880
rect 31937 8875 32003 8878
rect 38193 8875 38259 8878
rect 33777 8802 33843 8805
rect 34329 8802 34395 8805
rect 33777 8800 34395 8802
rect 33777 8744 33782 8800
rect 33838 8744 34334 8800
rect 34390 8744 34395 8800
rect 33777 8742 34395 8744
rect 33777 8739 33843 8742
rect 34329 8739 34395 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8530 800 8560
rect 2865 8530 2931 8533
rect 0 8528 2931 8530
rect 0 8472 2870 8528
rect 2926 8472 2931 8528
rect 0 8470 2931 8472
rect 0 8440 800 8470
rect 2865 8467 2931 8470
rect 32857 8530 32923 8533
rect 40033 8530 40099 8533
rect 32857 8528 40099 8530
rect 32857 8472 32862 8528
rect 32918 8472 40038 8528
rect 40094 8472 40099 8528
rect 32857 8470 40099 8472
rect 32857 8467 32923 8470
rect 40033 8467 40099 8470
rect 32029 8394 32095 8397
rect 35801 8394 35867 8397
rect 32029 8392 35867 8394
rect 32029 8336 32034 8392
rect 32090 8336 35806 8392
rect 35862 8336 35867 8392
rect 32029 8334 35867 8336
rect 32029 8331 32095 8334
rect 35801 8331 35867 8334
rect 37825 8394 37891 8397
rect 40953 8394 41019 8397
rect 37825 8392 41019 8394
rect 37825 8336 37830 8392
rect 37886 8336 40958 8392
rect 41014 8336 41019 8392
rect 37825 8334 41019 8336
rect 37825 8331 37891 8334
rect 40953 8331 41019 8334
rect 4208 8192 4528 8193
rect 0 8122 800 8152
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 21173 7850 21239 7853
rect 26877 7850 26943 7853
rect 21173 7848 26943 7850
rect 21173 7792 21178 7848
rect 21234 7792 26882 7848
rect 26938 7792 26943 7848
rect 21173 7790 26943 7792
rect 21173 7787 21239 7790
rect 26877 7787 26943 7790
rect 0 7714 800 7744
rect 1577 7714 1643 7717
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 0 7624 800 7654
rect 1577 7651 1643 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 0 7306 800 7336
rect 2957 7306 3023 7309
rect 0 7304 3023 7306
rect 0 7248 2962 7304
rect 3018 7248 3023 7304
rect 0 7246 3023 7248
rect 0 7216 800 7246
rect 2957 7243 3023 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 2313 6898 2379 6901
rect 0 6896 2379 6898
rect 0 6840 2318 6896
rect 2374 6840 2379 6896
rect 0 6838 2379 6840
rect 0 6808 800 6838
rect 2313 6835 2379 6838
rect 20989 6898 21055 6901
rect 22277 6898 22343 6901
rect 20989 6896 22343 6898
rect 20989 6840 20994 6896
rect 21050 6840 22282 6896
rect 22338 6840 22343 6896
rect 20989 6838 22343 6840
rect 20989 6835 21055 6838
rect 22277 6835 22343 6838
rect 38285 6626 38351 6629
rect 41689 6626 41755 6629
rect 38285 6624 41755 6626
rect 38285 6568 38290 6624
rect 38346 6568 41694 6624
rect 41750 6568 41755 6624
rect 38285 6566 41755 6568
rect 38285 6563 38351 6566
rect 41689 6563 41755 6566
rect 19568 6560 19888 6561
rect 0 6490 800 6520
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 1393 6490 1459 6493
rect 0 6488 1459 6490
rect 0 6432 1398 6488
rect 1454 6432 1459 6488
rect 0 6430 1459 6432
rect 0 6400 800 6430
rect 1393 6427 1459 6430
rect 30005 6490 30071 6493
rect 37365 6490 37431 6493
rect 30005 6488 37431 6490
rect 30005 6432 30010 6488
rect 30066 6432 37370 6488
rect 37426 6432 37431 6488
rect 30005 6430 37431 6432
rect 30005 6427 30071 6430
rect 37365 6427 37431 6430
rect 19885 6354 19951 6357
rect 27797 6354 27863 6357
rect 19885 6352 27863 6354
rect 19885 6296 19890 6352
rect 19946 6296 27802 6352
rect 27858 6296 27863 6352
rect 19885 6294 27863 6296
rect 19885 6291 19951 6294
rect 27797 6291 27863 6294
rect 29729 6218 29795 6221
rect 38561 6218 38627 6221
rect 29729 6216 38627 6218
rect 29729 6160 29734 6216
rect 29790 6160 38566 6216
rect 38622 6160 38627 6216
rect 29729 6158 38627 6160
rect 29729 6155 29795 6158
rect 38561 6155 38627 6158
rect 39389 6218 39455 6221
rect 47485 6218 47551 6221
rect 39389 6216 47551 6218
rect 39389 6160 39394 6216
rect 39450 6160 47490 6216
rect 47546 6160 47551 6216
rect 39389 6158 47551 6160
rect 39389 6155 39455 6158
rect 47485 6155 47551 6158
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 34697 5810 34763 5813
rect 35801 5810 35867 5813
rect 34697 5808 35867 5810
rect 34697 5752 34702 5808
rect 34758 5752 35806 5808
rect 35862 5752 35867 5808
rect 34697 5750 35867 5752
rect 34697 5747 34763 5750
rect 35801 5747 35867 5750
rect 41229 5810 41295 5813
rect 43345 5810 43411 5813
rect 41229 5808 43411 5810
rect 41229 5752 41234 5808
rect 41290 5752 43350 5808
rect 43406 5752 43411 5808
rect 41229 5750 43411 5752
rect 41229 5747 41295 5750
rect 43345 5747 43411 5750
rect 0 5674 800 5704
rect 1853 5674 1919 5677
rect 0 5672 1919 5674
rect 0 5616 1858 5672
rect 1914 5616 1919 5672
rect 0 5614 1919 5616
rect 0 5584 800 5614
rect 1853 5611 1919 5614
rect 24577 5674 24643 5677
rect 26969 5674 27035 5677
rect 24577 5672 27035 5674
rect 24577 5616 24582 5672
rect 24638 5616 26974 5672
rect 27030 5616 27035 5672
rect 24577 5614 27035 5616
rect 24577 5611 24643 5614
rect 26969 5611 27035 5614
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 0 5176 800 5296
rect 33593 5266 33659 5269
rect 36077 5266 36143 5269
rect 33593 5264 36143 5266
rect 33593 5208 33598 5264
rect 33654 5208 36082 5264
rect 36138 5208 36143 5264
rect 33593 5206 36143 5208
rect 33593 5203 33659 5206
rect 36077 5203 36143 5206
rect 23289 5130 23355 5133
rect 45737 5130 45803 5133
rect 23289 5128 45803 5130
rect 23289 5072 23294 5128
rect 23350 5072 45742 5128
rect 45798 5072 45803 5128
rect 23289 5070 45803 5072
rect 23289 5067 23355 5070
rect 45737 5067 45803 5070
rect 35341 4994 35407 4997
rect 36077 4994 36143 4997
rect 35341 4992 36143 4994
rect 35341 4936 35346 4992
rect 35402 4936 36082 4992
rect 36138 4936 36143 4992
rect 35341 4934 36143 4936
rect 35341 4931 35407 4934
rect 36077 4931 36143 4934
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 0 4722 800 4752
rect 2957 4722 3023 4725
rect 0 4720 3023 4722
rect 0 4664 2962 4720
rect 3018 4664 3023 4720
rect 0 4662 3023 4664
rect 0 4632 800 4662
rect 2957 4659 3023 4662
rect 35249 4722 35315 4725
rect 35709 4722 35775 4725
rect 35249 4720 35775 4722
rect 35249 4664 35254 4720
rect 35310 4664 35714 4720
rect 35770 4664 35775 4720
rect 35249 4662 35775 4664
rect 35249 4659 35315 4662
rect 35709 4659 35775 4662
rect 31109 4586 31175 4589
rect 33317 4586 33383 4589
rect 37733 4586 37799 4589
rect 31109 4584 37799 4586
rect 31109 4528 31114 4584
rect 31170 4528 33322 4584
rect 33378 4528 37738 4584
rect 37794 4528 37799 4584
rect 31109 4526 37799 4528
rect 31109 4523 31175 4526
rect 33317 4523 33383 4526
rect 37733 4523 37799 4526
rect 19568 4384 19888 4385
rect 0 4314 800 4344
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 2865 4314 2931 4317
rect 0 4312 2931 4314
rect 0 4256 2870 4312
rect 2926 4256 2931 4312
rect 0 4254 2931 4256
rect 0 4224 800 4254
rect 2865 4251 2931 4254
rect 3785 4178 3851 4181
rect 5533 4178 5599 4181
rect 3785 4176 5599 4178
rect 3785 4120 3790 4176
rect 3846 4120 5538 4176
rect 5594 4120 5599 4176
rect 3785 4118 5599 4120
rect 3785 4115 3851 4118
rect 5533 4115 5599 4118
rect 24669 4178 24735 4181
rect 38561 4178 38627 4181
rect 24669 4176 38627 4178
rect 24669 4120 24674 4176
rect 24730 4120 38566 4176
rect 38622 4120 38627 4176
rect 24669 4118 38627 4120
rect 24669 4115 24735 4118
rect 38561 4115 38627 4118
rect 40861 4178 40927 4181
rect 45829 4178 45895 4181
rect 46841 4178 46907 4181
rect 40861 4176 46907 4178
rect 40861 4120 40866 4176
rect 40922 4120 45834 4176
rect 45890 4120 46846 4176
rect 46902 4120 46907 4176
rect 40861 4118 46907 4120
rect 40861 4115 40927 4118
rect 45829 4115 45895 4118
rect 46841 4115 46907 4118
rect 22001 4042 22067 4045
rect 22185 4042 22251 4045
rect 22001 4040 22251 4042
rect 22001 3984 22006 4040
rect 22062 3984 22190 4040
rect 22246 3984 22251 4040
rect 22001 3982 22251 3984
rect 22001 3979 22067 3982
rect 22185 3979 22251 3982
rect 0 3906 800 3936
rect 1853 3906 1919 3909
rect 0 3904 1919 3906
rect 0 3848 1858 3904
rect 1914 3848 1919 3904
rect 0 3846 1919 3848
rect 0 3816 800 3846
rect 1853 3843 1919 3846
rect 20253 3906 20319 3909
rect 26969 3906 27035 3909
rect 20253 3904 27035 3906
rect 20253 3848 20258 3904
rect 20314 3848 26974 3904
rect 27030 3848 27035 3904
rect 20253 3846 27035 3848
rect 20253 3843 20319 3846
rect 26969 3843 27035 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 6913 3770 6979 3773
rect 12433 3770 12499 3773
rect 6913 3768 12499 3770
rect 6913 3712 6918 3768
rect 6974 3712 12438 3768
rect 12494 3712 12499 3768
rect 6913 3710 12499 3712
rect 6913 3707 6979 3710
rect 12433 3707 12499 3710
rect 22093 3770 22159 3773
rect 25405 3770 25471 3773
rect 22093 3768 25471 3770
rect 22093 3712 22098 3768
rect 22154 3712 25410 3768
rect 25466 3712 25471 3768
rect 22093 3710 25471 3712
rect 22093 3707 22159 3710
rect 25405 3707 25471 3710
rect 41321 3770 41387 3773
rect 42793 3770 42859 3773
rect 41321 3768 42859 3770
rect 41321 3712 41326 3768
rect 41382 3712 42798 3768
rect 42854 3712 42859 3768
rect 41321 3710 42859 3712
rect 41321 3707 41387 3710
rect 42793 3707 42859 3710
rect 43437 3770 43503 3773
rect 47577 3770 47643 3773
rect 43437 3768 47643 3770
rect 43437 3712 43442 3768
rect 43498 3712 47582 3768
rect 47638 3712 47643 3768
rect 43437 3710 47643 3712
rect 43437 3707 43503 3710
rect 47577 3707 47643 3710
rect 9213 3634 9279 3637
rect 10869 3634 10935 3637
rect 9213 3632 10935 3634
rect 9213 3576 9218 3632
rect 9274 3576 10874 3632
rect 10930 3576 10935 3632
rect 9213 3574 10935 3576
rect 9213 3571 9279 3574
rect 10869 3571 10935 3574
rect 22921 3634 22987 3637
rect 27981 3634 28047 3637
rect 22921 3632 28047 3634
rect 22921 3576 22926 3632
rect 22982 3576 27986 3632
rect 28042 3576 28047 3632
rect 22921 3574 28047 3576
rect 22921 3571 22987 3574
rect 27981 3571 28047 3574
rect 42149 3634 42215 3637
rect 47577 3634 47643 3637
rect 42149 3632 47643 3634
rect 42149 3576 42154 3632
rect 42210 3576 47582 3632
rect 47638 3576 47643 3632
rect 42149 3574 47643 3576
rect 42149 3571 42215 3574
rect 47577 3571 47643 3574
rect 48497 3634 48563 3637
rect 51165 3634 51231 3637
rect 48497 3632 51231 3634
rect 48497 3576 48502 3632
rect 48558 3576 51170 3632
rect 51226 3576 51231 3632
rect 48497 3574 51231 3576
rect 48497 3571 48563 3574
rect 51165 3571 51231 3574
rect 0 3408 800 3528
rect 2681 3498 2747 3501
rect 6453 3498 6519 3501
rect 2681 3496 6519 3498
rect 2681 3440 2686 3496
rect 2742 3440 6458 3496
rect 6514 3440 6519 3496
rect 2681 3438 6519 3440
rect 2681 3435 2747 3438
rect 6453 3435 6519 3438
rect 9121 3498 9187 3501
rect 10593 3498 10659 3501
rect 9121 3496 10659 3498
rect 9121 3440 9126 3496
rect 9182 3440 10598 3496
rect 10654 3440 10659 3496
rect 9121 3438 10659 3440
rect 9121 3435 9187 3438
rect 10593 3435 10659 3438
rect 45921 3498 45987 3501
rect 47209 3498 47275 3501
rect 47853 3498 47919 3501
rect 45921 3496 47919 3498
rect 45921 3440 45926 3496
rect 45982 3440 47214 3496
rect 47270 3440 47858 3496
rect 47914 3440 47919 3496
rect 45921 3438 47919 3440
rect 45921 3435 45987 3438
rect 47209 3435 47275 3438
rect 47853 3435 47919 3438
rect 48865 3498 48931 3501
rect 51533 3498 51599 3501
rect 48865 3496 51599 3498
rect 48865 3440 48870 3496
rect 48926 3440 51538 3496
rect 51594 3440 51599 3496
rect 48865 3438 51599 3440
rect 48865 3435 48931 3438
rect 51533 3435 51599 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 31017 3226 31083 3229
rect 36721 3226 36787 3229
rect 31017 3224 36787 3226
rect 31017 3168 31022 3224
rect 31078 3168 36726 3224
rect 36782 3168 36787 3224
rect 31017 3166 36787 3168
rect 31017 3163 31083 3166
rect 36721 3163 36787 3166
rect 39573 3226 39639 3229
rect 40861 3226 40927 3229
rect 42701 3226 42767 3229
rect 39573 3224 42767 3226
rect 39573 3168 39578 3224
rect 39634 3168 40866 3224
rect 40922 3168 42706 3224
rect 42762 3168 42767 3224
rect 39573 3166 42767 3168
rect 39573 3163 39639 3166
rect 40861 3163 40927 3166
rect 42701 3163 42767 3166
rect 0 3090 800 3120
rect 4061 3090 4127 3093
rect 0 3088 4127 3090
rect 0 3032 4066 3088
rect 4122 3032 4127 3088
rect 0 3030 4127 3032
rect 0 3000 800 3030
rect 4061 3027 4127 3030
rect 29821 3090 29887 3093
rect 31845 3090 31911 3093
rect 29821 3088 31911 3090
rect 29821 3032 29826 3088
rect 29882 3032 31850 3088
rect 31906 3032 31911 3088
rect 29821 3030 31911 3032
rect 29821 3027 29887 3030
rect 31845 3027 31911 3030
rect 35249 2954 35315 2957
rect 37917 2954 37983 2957
rect 35249 2952 37983 2954
rect 35249 2896 35254 2952
rect 35310 2896 37922 2952
rect 37978 2896 37983 2952
rect 35249 2894 37983 2896
rect 35249 2891 35315 2894
rect 37917 2891 37983 2894
rect 48773 2954 48839 2957
rect 55857 2954 55923 2957
rect 48773 2952 55923 2954
rect 48773 2896 48778 2952
rect 48834 2896 55862 2952
rect 55918 2896 55923 2952
rect 48773 2894 55923 2896
rect 48773 2891 48839 2894
rect 55857 2891 55923 2894
rect 4208 2752 4528 2753
rect 0 2682 800 2712
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 3693 2682 3759 2685
rect 0 2680 3759 2682
rect 0 2624 3698 2680
rect 3754 2624 3759 2680
rect 0 2622 3759 2624
rect 0 2592 800 2622
rect 3693 2619 3759 2622
rect 15193 2546 15259 2549
rect 19057 2546 19123 2549
rect 15193 2544 19123 2546
rect 15193 2488 15198 2544
rect 15254 2488 19062 2544
rect 19118 2488 19123 2544
rect 15193 2486 19123 2488
rect 15193 2483 15259 2486
rect 19057 2483 19123 2486
rect 10542 2348 10548 2412
rect 10612 2410 10618 2412
rect 51257 2410 51323 2413
rect 10612 2408 51323 2410
rect 10612 2352 51262 2408
rect 51318 2352 51323 2408
rect 10612 2350 51323 2352
rect 10612 2348 10618 2350
rect 51257 2347 51323 2350
rect 0 2274 800 2304
rect 3877 2274 3943 2277
rect 0 2272 3943 2274
rect 0 2216 3882 2272
rect 3938 2216 3943 2272
rect 0 2214 3943 2216
rect 0 2184 800 2214
rect 3877 2211 3943 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 0 1866 800 1896
rect 1853 1866 1919 1869
rect 0 1864 1919 1866
rect 0 1808 1858 1864
rect 1914 1808 1919 1864
rect 0 1806 1919 1808
rect 0 1776 800 1806
rect 1853 1803 1919 1806
rect 0 1458 800 1488
rect 3141 1458 3207 1461
rect 0 1456 3207 1458
rect 0 1400 3146 1456
rect 3202 1400 3207 1456
rect 0 1398 3207 1400
rect 0 1368 800 1398
rect 3141 1395 3207 1398
rect 0 1050 800 1080
rect 3325 1050 3391 1053
rect 0 1048 3391 1050
rect 0 992 3330 1048
rect 3386 992 3391 1048
rect 0 990 3391 992
rect 0 960 800 990
rect 3325 987 3391 990
rect 0 642 800 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 800 582
rect 1301 579 1367 582
rect 0 234 800 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 800 174
rect 2865 171 2931 174
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 10548 23488 10612 23492
rect 10548 23432 10562 23488
rect 10562 23432 10612 23488
rect 10548 23428 10612 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 9812 14512 9876 14516
rect 9812 14456 9826 14512
rect 9826 14456 9876 14512
rect 9812 14452 9876 14456
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 9812 12140 9876 12204
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 10548 2348 10612 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 19568 39200 19888 39760
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 10547 23492 10613 23493
rect 10547 23428 10548 23492
rect 10612 23428 10613 23492
rect 10547 23427 10613 23428
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 9811 14516 9877 14517
rect 9811 14452 9812 14516
rect 9876 14452 9877 14516
rect 9811 14451 9877 14452
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 9814 12205 9874 14451
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 10550 2413 10610 23427
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 10547 2412 10613 2413
rect 10547 2348 10548 2412
rect 10612 2348 10613 2412
rect 10547 2347 10613 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 39744 35248 39760
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 39200 50608 39760
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__fill_1  FILLER_0_3 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1644511149
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1644511149
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1644511149
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1644511149
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_236
timestamp 1644511149
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_244 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_347
timestamp 1644511149
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_355
timestamp 1644511149
transform 1 0 33764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1644511149
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1644511149
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1644511149
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1644511149
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1644511149
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1644511149
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1644511149
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1644511149
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_521
timestamp 1644511149
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1644511149
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_549
timestamp 1644511149
transform 1 0 51612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_567
timestamp 1644511149
transform 1 0 53268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_580
timestamp 1644511149
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_603
timestamp 1644511149
transform 1 0 56580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_611
timestamp 1644511149
transform 1 0 57316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1644511149
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1644511149
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1644511149
transform 1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1644511149
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_103
timestamp 1644511149
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_116
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_204
timestamp 1644511149
transform 1 0 19872 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1644511149
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1644511149
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_242
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_250
timestamp 1644511149
transform 1 0 24104 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_291 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_303
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_344
timestamp 1644511149
transform 1 0 32752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_350
timestamp 1644511149
transform 1 0 33304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1644511149
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1644511149
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_427
timestamp 1644511149
transform 1 0 40388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1644511149
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1644511149
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1644511149
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_481
timestamp 1644511149
transform 1 0 45356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1644511149
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_509
timestamp 1644511149
transform 1 0 47932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_521
timestamp 1644511149
transform 1 0 49036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_538
timestamp 1644511149
transform 1 0 50600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_546
timestamp 1644511149
transform 1 0 51336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_554
timestamp 1644511149
transform 1 0 52072 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_567
timestamp 1644511149
transform 1 0 53268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_583
timestamp 1644511149
transform 1 0 54740 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_599
timestamp 1644511149
transform 1 0 56212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_605
timestamp 1644511149
transform 1 0 56764 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_612
timestamp 1644511149
transform 1 0 57408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1644511149
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1644511149
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_33
timestamp 1644511149
transform 1 0 4140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_40
timestamp 1644511149
transform 1 0 4784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_47
timestamp 1644511149
transform 1 0 5428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_78
timestamp 1644511149
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_95
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1644511149
transform 1 0 15272 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_180
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_226
timestamp 1644511149
transform 1 0 21896 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1644511149
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_285
timestamp 1644511149
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_297
timestamp 1644511149
transform 1 0 28428 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1644511149
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_340
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_348
timestamp 1644511149
transform 1 0 33120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1644511149
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_390
timestamp 1644511149
transform 1 0 36984 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_402
timestamp 1644511149
transform 1 0 38088 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1644511149
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1644511149
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_427
timestamp 1644511149
transform 1 0 40388 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_432
timestamp 1644511149
transform 1 0 40848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_443
timestamp 1644511149
transform 1 0 41860 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1644511149
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_462
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1644511149
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_483
timestamp 1644511149
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1644511149
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_505
timestamp 1644511149
transform 1 0 47564 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_517
timestamp 1644511149
transform 1 0 48668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_549
timestamp 1644511149
transform 1 0 51612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_561
timestamp 1644511149
transform 1 0 52716 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_573
timestamp 1644511149
transform 1 0 53820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_585
timestamp 1644511149
transform 1 0 54924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1644511149
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_63
timestamp 1644511149
transform 1 0 6900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1644511149
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_82
timestamp 1644511149
transform 1 0 8648 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_95
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_121
timestamp 1644511149
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_129
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_142
timestamp 1644511149
transform 1 0 14168 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_153
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1644511149
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1644511149
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_209
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_221
timestamp 1644511149
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1644511149
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_248
timestamp 1644511149
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_260
timestamp 1644511149
transform 1 0 25024 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1644511149
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_343
timestamp 1644511149
transform 1 0 32660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_355
timestamp 1644511149
transform 1 0 33764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1644511149
transform 1 0 35972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_398
timestamp 1644511149
transform 1 0 37720 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_411
timestamp 1644511149
transform 1 0 38916 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_423
timestamp 1644511149
transform 1 0 40020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_431
timestamp 1644511149
transform 1 0 40756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_442
timestamp 1644511149
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_465
timestamp 1644511149
transform 1 0 43884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_477
timestamp 1644511149
transform 1 0 44988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_481
timestamp 1644511149
transform 1 0 45356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1644511149
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1644511149
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_525
timestamp 1644511149
transform 1 0 49404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_537
timestamp 1644511149
transform 1 0 50508 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_549
timestamp 1644511149
transform 1 0 51612 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_557
timestamp 1644511149
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1644511149
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1644511149
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_45
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1644511149
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_114
timestamp 1644511149
transform 1 0 11592 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_126
timestamp 1644511149
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1644511149
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_203
timestamp 1644511149
transform 1 0 19780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1644511149
transform 1 0 20884 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1644511149
transform 1 0 23092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_261
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_273
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_285
timestamp 1644511149
transform 1 0 27324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_293
timestamp 1644511149
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1644511149
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_322
timestamp 1644511149
transform 1 0 30728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_349
timestamp 1644511149
transform 1 0 33212 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_380
timestamp 1644511149
transform 1 0 36064 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_392
timestamp 1644511149
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1644511149
transform 1 0 37536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_428
timestamp 1644511149
transform 1 0 40480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_436
timestamp 1644511149
transform 1 0 41216 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_448
timestamp 1644511149
transform 1 0 42320 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_460
timestamp 1644511149
transform 1 0 43424 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1644511149
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_485
timestamp 1644511149
transform 1 0 45724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_507
timestamp 1644511149
transform 1 0 47748 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_515
timestamp 1644511149
transform 1 0 48484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_524
timestamp 1644511149
transform 1 0 49312 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1644511149
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_92
timestamp 1644511149
transform 1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1644511149
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1644511149
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_185
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_197
timestamp 1644511149
transform 1 0 19228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_203
timestamp 1644511149
transform 1 0 19780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_254
timestamp 1644511149
transform 1 0 24472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_265
timestamp 1644511149
transform 1 0 25484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1644511149
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_325
timestamp 1644511149
transform 1 0 31004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_355
timestamp 1644511149
transform 1 0 33764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_363
timestamp 1644511149
transform 1 0 34500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp 1644511149
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_426
timestamp 1644511149
transform 1 0 40296 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_438
timestamp 1644511149
transform 1 0 41400 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_446
timestamp 1644511149
transform 1 0 42136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_537
timestamp 1644511149
transform 1 0 50508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_556
timestamp 1644511149
transform 1 0 52256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_38
timestamp 1644511149
transform 1 0 4600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_50
timestamp 1644511149
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp 1644511149
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1644511149
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_102
timestamp 1644511149
transform 1 0 10488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_114
timestamp 1644511149
transform 1 0 11592 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_126
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1644511149
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1644511149
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1644511149
transform 1 0 16836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_183
timestamp 1644511149
transform 1 0 17940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_222
timestamp 1644511149
transform 1 0 21528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1644511149
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_241
timestamp 1644511149
transform 1 0 23276 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1644511149
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1644511149
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_325
timestamp 1644511149
transform 1 0 31004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_340
timestamp 1644511149
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_352
timestamp 1644511149
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_370
timestamp 1644511149
transform 1 0 35144 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_380
timestamp 1644511149
transform 1 0 36064 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_392
timestamp 1644511149
transform 1 0 37168 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_404
timestamp 1644511149
transform 1 0 38272 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_416
timestamp 1644511149
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_429
timestamp 1644511149
transform 1 0 40572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_440
timestamp 1644511149
transform 1 0 41584 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_460
timestamp 1644511149
transform 1 0 43424 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_472
timestamp 1644511149
transform 1 0 44528 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_482
timestamp 1644511149
transform 1 0 45448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_494
timestamp 1644511149
transform 1 0 46552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_504
timestamp 1644511149
transform 1 0 47472 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_516
timestamp 1644511149
transform 1 0 48576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_522
timestamp 1644511149
transform 1 0 49128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_530
timestamp 1644511149
transform 1 0 49864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_536
timestamp 1644511149
transform 1 0 50416 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_548
timestamp 1644511149
transform 1 0 51520 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_560
timestamp 1644511149
transform 1 0 52624 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_572
timestamp 1644511149
transform 1 0 53728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_584
timestamp 1644511149
transform 1 0 54832 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_14
timestamp 1644511149
transform 1 0 2392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_89
timestamp 1644511149
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1644511149
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_173
timestamp 1644511149
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1644511149
transform 1 0 18032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_196
timestamp 1644511149
transform 1 0 19136 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1644511149
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1644511149
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1644511149
transform 1 0 22448 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_244
timestamp 1644511149
transform 1 0 23552 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_256
timestamp 1644511149
transform 1 0 24656 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_268
timestamp 1644511149
transform 1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_274
timestamp 1644511149
transform 1 0 26312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_312
timestamp 1644511149
transform 1 0 29808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_320
timestamp 1644511149
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_357
timestamp 1644511149
transform 1 0 33948 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_364
timestamp 1644511149
transform 1 0 34592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_410
timestamp 1644511149
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_438
timestamp 1644511149
transform 1 0 41400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1644511149
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_462
timestamp 1644511149
transform 1 0 43608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_482
timestamp 1644511149
transform 1 0 45448 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_490
timestamp 1644511149
transform 1 0 46184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_499
timestamp 1644511149
transform 1 0 47012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_511
timestamp 1644511149
transform 1 0 48116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_534
timestamp 1644511149
transform 1 0 50232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_546
timestamp 1644511149
transform 1 0 51336 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_558
timestamp 1644511149
transform 1 0 52440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_13
timestamp 1644511149
transform 1 0 2300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_45
timestamp 1644511149
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1644511149
transform 1 0 6808 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1644511149
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1644511149
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1644511149
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1644511149
transform 1 0 12788 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1644511149
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_149
timestamp 1644511149
transform 1 0 14812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp 1644511149
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_183
timestamp 1644511149
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_212
timestamp 1644511149
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_224
timestamp 1644511149
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_231
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp 1644511149
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_341
timestamp 1644511149
transform 1 0 32476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_354
timestamp 1644511149
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1644511149
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_382
timestamp 1644511149
transform 1 0 36248 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_390
timestamp 1644511149
transform 1 0 36984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_396
timestamp 1644511149
transform 1 0 37536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_405
timestamp 1644511149
transform 1 0 38364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1644511149
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_444
timestamp 1644511149
transform 1 0 41952 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_493
timestamp 1644511149
transform 1 0 46460 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_510
timestamp 1644511149
transform 1 0 48024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_518
timestamp 1644511149
transform 1 0 48760 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_523
timestamp 1644511149
transform 1 0 49220 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_536
timestamp 1644511149
transform 1 0 50416 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_544
timestamp 1644511149
transform 1 0 51152 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_561
timestamp 1644511149
transform 1 0 52716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_573
timestamp 1644511149
transform 1 0 53820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_585
timestamp 1644511149
transform 1 0 54924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1644511149
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_21
timestamp 1644511149
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_33
timestamp 1644511149
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1644511149
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_73
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_85
timestamp 1644511149
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1644511149
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_144
timestamp 1644511149
transform 1 0 14352 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1644511149
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_201
timestamp 1644511149
transform 1 0 19596 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1644511149
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1644511149
transform 1 0 22356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_242
timestamp 1644511149
transform 1 0 23368 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_263
timestamp 1644511149
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1644511149
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_298
timestamp 1644511149
transform 1 0 28520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_310
timestamp 1644511149
transform 1 0 29624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_322
timestamp 1644511149
transform 1 0 30728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1644511149
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_345
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_351
timestamp 1644511149
transform 1 0 33396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_356
timestamp 1644511149
transform 1 0 33856 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_368
timestamp 1644511149
transform 1 0 34960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_372
timestamp 1644511149
transform 1 0 35328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_375
timestamp 1644511149
transform 1 0 35604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1644511149
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1644511149
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_401
timestamp 1644511149
transform 1 0 37996 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_411
timestamp 1644511149
transform 1 0 38916 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_423
timestamp 1644511149
transform 1 0 40020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_435
timestamp 1644511149
transform 1 0 41124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_479
timestamp 1644511149
transform 1 0 45172 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_487
timestamp 1644511149
transform 1 0 45908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_496
timestamp 1644511149
transform 1 0 46736 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_567
timestamp 1644511149
transform 1 0 53268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_579
timestamp 1644511149
transform 1 0 54372 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_591
timestamp 1644511149
transform 1 0 55476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_603
timestamp 1644511149
transform 1 0 56580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_35
timestamp 1644511149
transform 1 0 4324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_47
timestamp 1644511149
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_100
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_110
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_119
timestamp 1644511149
transform 1 0 12052 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1644511149
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_151
timestamp 1644511149
transform 1 0 14996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1644511149
transform 1 0 16100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1644511149
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1644511149
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1644511149
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_217
timestamp 1644511149
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_226
timestamp 1644511149
transform 1 0 21896 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_238
timestamp 1644511149
transform 1 0 23000 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1644511149
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1644511149
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_274
timestamp 1644511149
transform 1 0 26312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_284
timestamp 1644511149
transform 1 0 27232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_295
timestamp 1644511149
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1644511149
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1644511149
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_381
timestamp 1644511149
transform 1 0 36156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_386
timestamp 1644511149
transform 1 0 36616 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1644511149
transform 1 0 37720 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_410
timestamp 1644511149
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1644511149
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_456
timestamp 1644511149
transform 1 0 43056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_468
timestamp 1644511149
transform 1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_539
timestamp 1644511149
transform 1 0 50692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_551
timestamp 1644511149
transform 1 0 51796 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_559
timestamp 1644511149
transform 1 0 52532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_576
timestamp 1644511149
transform 1 0 54096 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_12
timestamp 1644511149
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1644511149
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1644511149
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_85
timestamp 1644511149
transform 1 0 8924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1644511149
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1644511149
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_138
timestamp 1644511149
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_176
timestamp 1644511149
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_188
timestamp 1644511149
transform 1 0 18400 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_200
timestamp 1644511149
transform 1 0 19504 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_212
timestamp 1644511149
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1644511149
transform 1 0 23460 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_248
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_260
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1644511149
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_285
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_289
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1644511149
transform 1 0 28520 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1644511149
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_327
timestamp 1644511149
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_355
timestamp 1644511149
transform 1 0 33764 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_372
timestamp 1644511149
transform 1 0 35328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_396
timestamp 1644511149
transform 1 0 37536 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_404
timestamp 1644511149
transform 1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_416
timestamp 1644511149
transform 1 0 39376 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_430
timestamp 1644511149
transform 1 0 40664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_442
timestamp 1644511149
transform 1 0 41768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_458
timestamp 1644511149
transform 1 0 43240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_470
timestamp 1644511149
transform 1 0 44344 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_498
timestamp 1644511149
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_523
timestamp 1644511149
transform 1 0 49220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_540
timestamp 1644511149
transform 1 0 50784 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_552
timestamp 1644511149
transform 1 0 51888 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_570
timestamp 1644511149
transform 1 0 53544 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_582
timestamp 1644511149
transform 1 0 54648 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_594
timestamp 1644511149
transform 1 0 55752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_606
timestamp 1644511149
transform 1 0 56856 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1644511149
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1644511149
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_35
timestamp 1644511149
transform 1 0 4324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_47
timestamp 1644511149
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_59
timestamp 1644511149
transform 1 0 6532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_63
timestamp 1644511149
transform 1 0 6900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1644511149
transform 1 0 7544 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1644511149
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1644511149
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_108
timestamp 1644511149
transform 1 0 11040 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_120
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1644511149
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_148
timestamp 1644511149
transform 1 0 14720 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1644511149
transform 1 0 15824 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_175
timestamp 1644511149
transform 1 0 17204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_205
timestamp 1644511149
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_214
timestamp 1644511149
transform 1 0 20792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_241
timestamp 1644511149
transform 1 0 23276 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_261
timestamp 1644511149
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1644511149
transform 1 0 27048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1644511149
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1644511149
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_330
timestamp 1644511149
transform 1 0 31464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_343
timestamp 1644511149
transform 1 0 32660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_355
timestamp 1644511149
transform 1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1644511149
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_375
timestamp 1644511149
transform 1 0 35604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1644511149
transform 1 0 36524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_397
timestamp 1644511149
transform 1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1644511149
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_441
timestamp 1644511149
transform 1 0 41676 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_451
timestamp 1644511149
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_463
timestamp 1644511149
transform 1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_480
timestamp 1644511149
transform 1 0 45264 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_492
timestamp 1644511149
transform 1 0 46368 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_504
timestamp 1644511149
transform 1 0 47472 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_516
timestamp 1644511149
transform 1 0 48576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1644511149
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_537
timestamp 1644511149
transform 1 0 50508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_549
timestamp 1644511149
transform 1 0 51612 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_558
timestamp 1644511149
transform 1 0 52440 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_570
timestamp 1644511149
transform 1 0 53544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_576
timestamp 1644511149
transform 1 0 54096 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_19
timestamp 1644511149
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1644511149
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_63
timestamp 1644511149
transform 1 0 6900 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1644511149
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_83
timestamp 1644511149
transform 1 0 8740 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_87
timestamp 1644511149
transform 1 0 9108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1644511149
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_121
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1644511149
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_153
timestamp 1644511149
transform 1 0 15180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1644511149
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1644511149
transform 1 0 17572 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_196
timestamp 1644511149
transform 1 0 19136 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1644511149
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_244
timestamp 1644511149
transform 1 0 23552 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_256
timestamp 1644511149
transform 1 0 24656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_310
timestamp 1644511149
transform 1 0 29624 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_318
timestamp 1644511149
transform 1 0 30360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_326
timestamp 1644511149
transform 1 0 31096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1644511149
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_343
timestamp 1644511149
transform 1 0 32660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_346
timestamp 1644511149
transform 1 0 32936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_355
timestamp 1644511149
transform 1 0 33764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_364
timestamp 1644511149
transform 1 0 34592 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_372
timestamp 1644511149
transform 1 0 35328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1644511149
transform 1 0 35972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_399
timestamp 1644511149
transform 1 0 37812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_407
timestamp 1644511149
transform 1 0 38548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_416
timestamp 1644511149
transform 1 0 39376 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_428
timestamp 1644511149
transform 1 0 40480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_432
timestamp 1644511149
transform 1 0 40848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_440
timestamp 1644511149
transform 1 0 41584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_454
timestamp 1644511149
transform 1 0 42872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_466
timestamp 1644511149
transform 1 0 43976 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_478
timestamp 1644511149
transform 1 0 45080 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_486
timestamp 1644511149
transform 1 0 45816 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_498
timestamp 1644511149
transform 1 0 46920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_513
timestamp 1644511149
transform 1 0 48300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_520
timestamp 1644511149
transform 1 0 48944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_530
timestamp 1644511149
transform 1 0 49864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_542
timestamp 1644511149
transform 1 0 50968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_551
timestamp 1644511149
transform 1 0 51796 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_564
timestamp 1644511149
transform 1 0 52992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_577
timestamp 1644511149
transform 1 0 54188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_581
timestamp 1644511149
transform 1 0 54556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_601
timestamp 1644511149
transform 1 0 56396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_613
timestamp 1644511149
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1644511149
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_37
timestamp 1644511149
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_56
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_67
timestamp 1644511149
transform 1 0 7268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1644511149
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_120
timestamp 1644511149
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1644511149
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1644511149
transform 1 0 15272 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_166
timestamp 1644511149
transform 1 0 16376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_174
timestamp 1644511149
transform 1 0 17112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_179
timestamp 1644511149
transform 1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_275
timestamp 1644511149
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_287
timestamp 1644511149
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1644511149
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_344
timestamp 1644511149
transform 1 0 32752 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_356
timestamp 1644511149
transform 1 0 33856 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_369
timestamp 1644511149
transform 1 0 35052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_375
timestamp 1644511149
transform 1 0 35604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_383
timestamp 1644511149
transform 1 0 36340 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_395
timestamp 1644511149
transform 1 0 37444 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_408
timestamp 1644511149
transform 1 0 38640 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_440
timestamp 1644511149
transform 1 0 41584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_449
timestamp 1644511149
transform 1 0 42412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_471
timestamp 1644511149
transform 1 0 44436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_483
timestamp 1644511149
transform 1 0 45540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_508
timestamp 1644511149
transform 1 0 47840 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_520
timestamp 1644511149
transform 1 0 48944 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1644511149
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1644511149
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1644511149
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_71
timestamp 1644511149
transform 1 0 7636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_79
timestamp 1644511149
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_91
timestamp 1644511149
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_103
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1644511149
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1644511149
transform 1 0 13524 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_195
timestamp 1644511149
transform 1 0 19044 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1644511149
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1644511149
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_323
timestamp 1644511149
transform 1 0 30820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_331
timestamp 1644511149
transform 1 0 31556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_377
timestamp 1644511149
transform 1 0 35788 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1644511149
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_455
timestamp 1644511149
transform 1 0 42964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_467
timestamp 1644511149
transform 1 0 44068 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_479
timestamp 1644511149
transform 1 0 45172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_491
timestamp 1644511149
transform 1 0 46276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_526
timestamp 1644511149
transform 1 0 49496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_535
timestamp 1644511149
transform 1 0 50324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_547
timestamp 1644511149
transform 1 0 51428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_580
timestamp 1644511149
transform 1 0 54464 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_592
timestamp 1644511149
transform 1 0 55568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_604
timestamp 1644511149
transform 1 0 56672 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1644511149
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1644511149
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1644511149
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_158
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_167
timestamp 1644511149
transform 1 0 16468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1644511149
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1644511149
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1644511149
transform 1 0 20700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1644511149
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_234
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_258
timestamp 1644511149
transform 1 0 24840 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_267
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1644511149
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1644511149
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_325
timestamp 1644511149
transform 1 0 31004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_342
timestamp 1644511149
transform 1 0 32568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_353
timestamp 1644511149
transform 1 0 33580 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1644511149
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_369
timestamp 1644511149
transform 1 0 35052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_376
timestamp 1644511149
transform 1 0 35696 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_387
timestamp 1644511149
transform 1 0 36708 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_399
timestamp 1644511149
transform 1 0 37812 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_411
timestamp 1644511149
transform 1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_438
timestamp 1644511149
transform 1 0 41400 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_450
timestamp 1644511149
transform 1 0 42504 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_462
timestamp 1644511149
transform 1 0 43608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1644511149
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_508
timestamp 1644511149
transform 1 0 47840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_528
timestamp 1644511149
transform 1 0 49680 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_544
timestamp 1644511149
transform 1 0 51152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_556
timestamp 1644511149
transform 1 0 52256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_568
timestamp 1644511149
transform 1 0 53360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_572
timestamp 1644511149
transform 1 0 53728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_584
timestamp 1644511149
transform 1 0 54832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_6
timestamp 1644511149
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_14
timestamp 1644511149
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1644511149
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1644511149
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_63
timestamp 1644511149
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_72
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_76
timestamp 1644511149
transform 1 0 8096 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_85
timestamp 1644511149
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1644511149
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1644511149
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1644511149
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_121
timestamp 1644511149
transform 1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_141
timestamp 1644511149
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_182
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_208
timestamp 1644511149
transform 1 0 20240 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1644511149
transform 1 0 23276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_253
timestamp 1644511149
transform 1 0 24380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1644511149
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_288
timestamp 1644511149
transform 1 0 27600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_296
timestamp 1644511149
transform 1 0 28336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_308
timestamp 1644511149
transform 1 0 29440 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_318
timestamp 1644511149
transform 1 0 30360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1644511149
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_341
timestamp 1644511149
transform 1 0 32476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_353
timestamp 1644511149
transform 1 0 33580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_362
timestamp 1644511149
transform 1 0 34408 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_382
timestamp 1644511149
transform 1 0 36248 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1644511149
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_398
timestamp 1644511149
transform 1 0 37720 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_409
timestamp 1644511149
transform 1 0 38732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_418
timestamp 1644511149
transform 1 0 39560 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_424
timestamp 1644511149
transform 1 0 40112 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_431
timestamp 1644511149
transform 1 0 40756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1644511149
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_465
timestamp 1644511149
transform 1 0 43884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_479
timestamp 1644511149
transform 1 0 45172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_491
timestamp 1644511149
transform 1 0 46276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_518
timestamp 1644511149
transform 1 0 48760 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_530
timestamp 1644511149
transform 1 0 49864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_542
timestamp 1644511149
transform 1 0 50968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_546
timestamp 1644511149
transform 1 0 51336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_552
timestamp 1644511149
transform 1 0 51888 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_567
timestamp 1644511149
transform 1 0 53268 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_570
timestamp 1644511149
transform 1 0 53544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_577
timestamp 1644511149
transform 1 0 54188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_591
timestamp 1644511149
transform 1 0 55476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1644511149
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_12
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp 1644511149
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_37
timestamp 1644511149
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_45
timestamp 1644511149
transform 1 0 5244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_56
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1644511149
transform 1 0 6992 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_70
timestamp 1644511149
transform 1 0 7544 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_91
timestamp 1644511149
transform 1 0 9476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_103
timestamp 1644511149
transform 1 0 10580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_161
timestamp 1644511149
transform 1 0 15916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_173
timestamp 1644511149
transform 1 0 17020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_181
timestamp 1644511149
transform 1 0 17756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_225
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_231
timestamp 1644511149
transform 1 0 22356 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1644511149
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_269
timestamp 1644511149
transform 1 0 25852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_278
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_286
timestamp 1644511149
transform 1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_291
timestamp 1644511149
transform 1 0 27876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1644511149
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_329
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_334
timestamp 1644511149
transform 1 0 31832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_344
timestamp 1644511149
transform 1 0 32752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_348
timestamp 1644511149
transform 1 0 33120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_356
timestamp 1644511149
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_380
timestamp 1644511149
transform 1 0 36064 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_391
timestamp 1644511149
transform 1 0 37076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1644511149
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_425
timestamp 1644511149
transform 1 0 40204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_464
timestamp 1644511149
transform 1 0 43792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_472
timestamp 1644511149
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_496
timestamp 1644511149
transform 1 0 46736 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_508
timestamp 1644511149
transform 1 0 47840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_516
timestamp 1644511149
transform 1 0 48576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_522
timestamp 1644511149
transform 1 0 49128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_530
timestamp 1644511149
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_539
timestamp 1644511149
transform 1 0 50692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_554
timestamp 1644511149
transform 1 0 52072 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_566
timestamp 1644511149
transform 1 0 53176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_577
timestamp 1644511149
transform 1 0 54188 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_585
timestamp 1644511149
transform 1 0 54924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_593
timestamp 1644511149
transform 1 0 55660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_605
timestamp 1644511149
transform 1 0 56764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_617
timestamp 1644511149
transform 1 0 57868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_18
timestamp 1644511149
transform 1 0 2760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_74
timestamp 1644511149
transform 1 0 7912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_88
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_94
timestamp 1644511149
transform 1 0 9752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1644511149
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1644511149
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_126
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_139
timestamp 1644511149
transform 1 0 13892 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_147
timestamp 1644511149
transform 1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1644511149
transform 1 0 15088 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1644511149
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1644511149
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_254
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_266
timestamp 1644511149
transform 1 0 25576 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1644511149
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_301
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_313
timestamp 1644511149
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1644511149
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1644511149
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_412
timestamp 1644511149
transform 1 0 39008 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_425
timestamp 1644511149
transform 1 0 40204 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_443
timestamp 1644511149
transform 1 0 41860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_474
timestamp 1644511149
transform 1 0 44712 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_480
timestamp 1644511149
transform 1 0 45264 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_484
timestamp 1644511149
transform 1 0 45632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_496
timestamp 1644511149
transform 1 0 46736 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_514
timestamp 1644511149
transform 1 0 48392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_534
timestamp 1644511149
transform 1 0 50232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_543
timestamp 1644511149
transform 1 0 51060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_555
timestamp 1644511149
transform 1 0 52164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_569
timestamp 1644511149
transform 1 0 53452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_575
timestamp 1644511149
transform 1 0 54004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_581
timestamp 1644511149
transform 1 0 54556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_586
timestamp 1644511149
transform 1 0 55016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_594
timestamp 1644511149
transform 1 0 55752 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_611
timestamp 1644511149
transform 1 0 57316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp 1644511149
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_45
timestamp 1644511149
transform 1 0 5244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_57
timestamp 1644511149
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1644511149
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_103
timestamp 1644511149
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_110
timestamp 1644511149
transform 1 0 11224 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_122
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1644511149
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_145
timestamp 1644511149
transform 1 0 14444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_169
timestamp 1644511149
transform 1 0 16652 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_175
timestamp 1644511149
transform 1 0 17204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_212
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_218
timestamp 1644511149
transform 1 0 21160 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_261
timestamp 1644511149
transform 1 0 25116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_285
timestamp 1644511149
transform 1 0 27324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_296
timestamp 1644511149
transform 1 0 28336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_317
timestamp 1644511149
transform 1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_325
timestamp 1644511149
transform 1 0 31004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_341
timestamp 1644511149
transform 1 0 32476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1644511149
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_375
timestamp 1644511149
transform 1 0 35604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_388
timestamp 1644511149
transform 1 0 36800 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_400
timestamp 1644511149
transform 1 0 37904 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1644511149
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_428
timestamp 1644511149
transform 1 0 40480 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_434
timestamp 1644511149
transform 1 0 41032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_451
timestamp 1644511149
transform 1 0 42596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_463
timestamp 1644511149
transform 1 0 43700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1644511149
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_493
timestamp 1644511149
transform 1 0 46460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_505
timestamp 1644511149
transform 1 0 47564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_517
timestamp 1644511149
transform 1 0 48668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_521
timestamp 1644511149
transform 1 0 49036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_538
timestamp 1644511149
transform 1 0 50600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_550
timestamp 1644511149
transform 1 0 51704 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_562
timestamp 1644511149
transform 1 0 52808 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_575
timestamp 1644511149
transform 1 0 54004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_583
timestamp 1644511149
transform 1 0 54740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_14
timestamp 1644511149
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_88
timestamp 1644511149
transform 1 0 9200 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_100
timestamp 1644511149
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1644511149
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1644511149
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1644511149
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1644511149
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_341
timestamp 1644511149
transform 1 0 32476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1644511149
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_379
timestamp 1644511149
transform 1 0 35972 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1644511149
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_427
timestamp 1644511149
transform 1 0 40388 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_435
timestamp 1644511149
transform 1 0 41124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_477
timestamp 1644511149
transform 1 0 44988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_483
timestamp 1644511149
transform 1 0 45540 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_489
timestamp 1644511149
transform 1 0 46092 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1644511149
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_540
timestamp 1644511149
transform 1 0 50784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_552
timestamp 1644511149
transform 1 0 51888 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_565
timestamp 1644511149
transform 1 0 53084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_582
timestamp 1644511149
transform 1 0 54648 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_594
timestamp 1644511149
transform 1 0 55752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_606
timestamp 1644511149
transform 1 0 56856 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_614
timestamp 1644511149
transform 1 0 57592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1644511149
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_50
timestamp 1644511149
transform 1 0 5704 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_62
timestamp 1644511149
transform 1 0 6808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1644511149
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1644511149
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1644511149
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_130
timestamp 1644511149
transform 1 0 13064 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_169
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_241
timestamp 1644511149
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp 1644511149
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1644511149
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_275
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1644511149
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1644511149
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_336
timestamp 1644511149
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_348
timestamp 1644511149
transform 1 0 33120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1644511149
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_386
timestamp 1644511149
transform 1 0 36616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_397
timestamp 1644511149
transform 1 0 37628 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_409
timestamp 1644511149
transform 1 0 38732 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_417
timestamp 1644511149
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_430
timestamp 1644511149
transform 1 0 40664 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_442
timestamp 1644511149
transform 1 0 41768 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_454
timestamp 1644511149
transform 1 0 42872 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_466
timestamp 1644511149
transform 1 0 43976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1644511149
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_493
timestamp 1644511149
transform 1 0 46460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_510
timestamp 1644511149
transform 1 0 48024 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_522
timestamp 1644511149
transform 1 0 49128 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_530
timestamp 1644511149
transform 1 0 49864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_549
timestamp 1644511149
transform 1 0 51612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_561
timestamp 1644511149
transform 1 0 52716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_574
timestamp 1644511149
transform 1 0 53912 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_586
timestamp 1644511149
transform 1 0 55016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_25
timestamp 1644511149
transform 1 0 3404 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_33
timestamp 1644511149
transform 1 0 4140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1644511149
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1644511149
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1644511149
transform 1 0 9016 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1644511149
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1644511149
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_121
timestamp 1644511149
transform 1 0 12236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_128
timestamp 1644511149
transform 1 0 12880 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_140
timestamp 1644511149
transform 1 0 13984 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_146
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1644511149
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_234
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_262
timestamp 1644511149
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_296
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_308
timestamp 1644511149
transform 1 0 29440 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_320
timestamp 1644511149
transform 1 0 30544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1644511149
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_366
timestamp 1644511149
transform 1 0 34776 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_378
timestamp 1644511149
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1644511149
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_410
timestamp 1644511149
transform 1 0 38824 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_422
timestamp 1644511149
transform 1 0 39928 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_430
timestamp 1644511149
transform 1 0 40664 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_435
timestamp 1644511149
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_457
timestamp 1644511149
transform 1 0 43148 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_463
timestamp 1644511149
transform 1 0 43700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_471
timestamp 1644511149
transform 1 0 44436 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_483
timestamp 1644511149
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_495
timestamp 1644511149
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_520
timestamp 1644511149
transform 1 0 48944 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_532
timestamp 1644511149
transform 1 0 50048 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_544
timestamp 1644511149
transform 1 0 51152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_556
timestamp 1644511149
transform 1 0 52256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_567
timestamp 1644511149
transform 1 0 53268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_579
timestamp 1644511149
transform 1 0 54372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_591
timestamp 1644511149
transform 1 0 55476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_603
timestamp 1644511149
transform 1 0 56580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1644511149
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1644511149
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1644511149
transform 1 0 6808 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_74
timestamp 1644511149
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1644511149
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1644511149
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1644511149
transform 1 0 15548 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1644511149
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_178
timestamp 1644511149
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_184
timestamp 1644511149
transform 1 0 18032 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_204
timestamp 1644511149
transform 1 0 19872 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_216
timestamp 1644511149
transform 1 0 20976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_224
timestamp 1644511149
transform 1 0 21712 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_231
timestamp 1644511149
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_272
timestamp 1644511149
transform 1 0 26128 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_279
timestamp 1644511149
transform 1 0 26772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_288
timestamp 1644511149
transform 1 0 27600 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1644511149
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_319
timestamp 1644511149
transform 1 0 30452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_331
timestamp 1644511149
transform 1 0 31556 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_343
timestamp 1644511149
transform 1 0 32660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_351
timestamp 1644511149
transform 1 0 33396 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1644511149
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_371
timestamp 1644511149
transform 1 0 35236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_375
timestamp 1644511149
transform 1 0 35604 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_386
timestamp 1644511149
transform 1 0 36616 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_394
timestamp 1644511149
transform 1 0 37352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_430
timestamp 1644511149
transform 1 0 40664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_449
timestamp 1644511149
transform 1 0 42412 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_464
timestamp 1644511149
transform 1 0 43792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_565
timestamp 1644511149
transform 1 0 53084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_584
timestamp 1644511149
transform 1 0 54832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_23
timestamp 1644511149
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_35
timestamp 1644511149
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1644511149
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_73
timestamp 1644511149
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_85
timestamp 1644511149
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_97
timestamp 1644511149
transform 1 0 10028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_136
timestamp 1644511149
transform 1 0 13616 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191
timestamp 1644511149
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1644511149
transform 1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_241
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_264
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_302
timestamp 1644511149
transform 1 0 28888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_322
timestamp 1644511149
transform 1 0 30728 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_344
timestamp 1644511149
transform 1 0 32752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1644511149
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_375
timestamp 1644511149
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 1644511149
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_425
timestamp 1644511149
transform 1 0 40204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_442
timestamp 1644511149
transform 1 0 41768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_468
timestamp 1644511149
transform 1 0 44160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_477
timestamp 1644511149
transform 1 0 44988 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_489
timestamp 1644511149
transform 1 0 46092 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_493
timestamp 1644511149
transform 1 0 46460 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_500
timestamp 1644511149
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_512
timestamp 1644511149
transform 1 0 48208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_91
timestamp 1644511149
transform 1 0 9476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_103
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_122
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1644511149
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_173
timestamp 1644511149
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_314
timestamp 1644511149
transform 1 0 29992 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_325
timestamp 1644511149
transform 1 0 31004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1644511149
transform 1 0 32108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_349
timestamp 1644511149
transform 1 0 33212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1644511149
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_375
timestamp 1644511149
transform 1 0 35604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_379
timestamp 1644511149
transform 1 0 35972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_394
timestamp 1644511149
transform 1 0 37352 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_406
timestamp 1644511149
transform 1 0 38456 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1644511149
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_429
timestamp 1644511149
transform 1 0 40572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_436
timestamp 1644511149
transform 1 0 41216 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_448
timestamp 1644511149
transform 1 0 42320 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_468
timestamp 1644511149
transform 1 0 44160 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_484
timestamp 1644511149
transform 1 0 45632 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_492
timestamp 1644511149
transform 1 0 46368 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_502
timestamp 1644511149
transform 1 0 47288 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_508
timestamp 1644511149
transform 1 0 47840 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_524
timestamp 1644511149
transform 1 0 49312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_18
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_88
timestamp 1644511149
transform 1 0 9200 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_100
timestamp 1644511149
transform 1 0 10304 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_124
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1644511149
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_147
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_153
timestamp 1644511149
transform 1 0 15180 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1644511149
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_201
timestamp 1644511149
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1644511149
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_233
timestamp 1644511149
transform 1 0 22540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_253
timestamp 1644511149
transform 1 0 24380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_264
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_301
timestamp 1644511149
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_313
timestamp 1644511149
transform 1 0 29900 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_321
timestamp 1644511149
transform 1 0 30636 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_345
timestamp 1644511149
transform 1 0 32844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_357
timestamp 1644511149
transform 1 0 33948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_369
timestamp 1644511149
transform 1 0 35052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1644511149
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1644511149
transform 1 0 39008 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1644511149
transform 1 0 40112 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1644511149
transform 1 0 41216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_453
timestamp 1644511149
transform 1 0 42780 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_457
timestamp 1644511149
transform 1 0 43148 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_469
timestamp 1644511149
transform 1 0 44252 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_477
timestamp 1644511149
transform 1 0 44988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_483
timestamp 1644511149
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_495
timestamp 1644511149
transform 1 0 46644 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_13
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1644511149
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1644511149
transform 1 0 4048 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1644511149
transform 1 0 6256 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_91
timestamp 1644511149
transform 1 0 9476 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_103
timestamp 1644511149
transform 1 0 10580 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_115
timestamp 1644511149
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_119
timestamp 1644511149
transform 1 0 12052 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1644511149
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_182
timestamp 1644511149
transform 1 0 17848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_207
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1644511149
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1644511149
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1644511149
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_314
timestamp 1644511149
transform 1 0 29992 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_326
timestamp 1644511149
transform 1 0 31096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_334
timestamp 1644511149
transform 1 0 31832 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_346
timestamp 1644511149
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_369
timestamp 1644511149
transform 1 0 35052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_397
timestamp 1644511149
transform 1 0 37628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_409
timestamp 1644511149
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_417
timestamp 1644511149
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_427
timestamp 1644511149
transform 1 0 40388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_439
timestamp 1644511149
transform 1 0 41492 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_467
timestamp 1644511149
transform 1 0 44068 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_481
timestamp 1644511149
transform 1 0 45356 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_498
timestamp 1644511149
transform 1 0 46920 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_510
timestamp 1644511149
transform 1 0 48024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_517
timestamp 1644511149
transform 1 0 48668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_529
timestamp 1644511149
transform 1 0 49772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1644511149
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_67
timestamp 1644511149
transform 1 0 7268 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_75
timestamp 1644511149
transform 1 0 8004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_119
timestamp 1644511149
transform 1 0 12052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_131
timestamp 1644511149
transform 1 0 13156 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_143
timestamp 1644511149
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_298
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_302
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_307
timestamp 1644511149
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_319
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_323
timestamp 1644511149
transform 1 0 30820 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_363
timestamp 1644511149
transform 1 0 34500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_377
timestamp 1644511149
transform 1 0 35788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1644511149
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_396
timestamp 1644511149
transform 1 0 37536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_408
timestamp 1644511149
transform 1 0 38640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_413
timestamp 1644511149
transform 1 0 39100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_424
timestamp 1644511149
transform 1 0 40112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_444
timestamp 1644511149
transform 1 0 41952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1644511149
transform 1 0 6716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1644511149
transform 1 0 7452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1644511149
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_88
timestamp 1644511149
transform 1 0 9200 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_103
timestamp 1644511149
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1644511149
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_128
timestamp 1644511149
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_162
timestamp 1644511149
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_174
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1644511149
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1644511149
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_218
timestamp 1644511149
transform 1 0 21160 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_226
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_235
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1644511149
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_317
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_329
timestamp 1644511149
transform 1 0 31372 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 1644511149
transform 1 0 31924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_344
timestamp 1644511149
transform 1 0 32752 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1644511149
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_375
timestamp 1644511149
transform 1 0 35604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_388
timestamp 1644511149
transform 1 0 36800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_428
timestamp 1644511149
transform 1 0 40480 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_440
timestamp 1644511149
transform 1 0 41584 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_452
timestamp 1644511149
transform 1 0 42688 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_464
timestamp 1644511149
transform 1 0 43792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_6
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_21
timestamp 1644511149
transform 1 0 3036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_33
timestamp 1644511149
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1644511149
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_67
timestamp 1644511149
transform 1 0 7268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_77
timestamp 1644511149
transform 1 0 8188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1644511149
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_141
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_177
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1644511149
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1644511149
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1644511149
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_253
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_262
timestamp 1644511149
transform 1 0 25208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_266
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_269
timestamp 1644511149
transform 1 0 25852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_290
timestamp 1644511149
transform 1 0 27784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_302
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_311
timestamp 1644511149
transform 1 0 29716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_321
timestamp 1644511149
transform 1 0 30636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1644511149
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_359
timestamp 1644511149
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_381
timestamp 1644511149
transform 1 0 36156 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_415
timestamp 1644511149
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_427
timestamp 1644511149
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1644511149
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1644511149
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1644511149
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_45
timestamp 1644511149
transform 1 0 5244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_117
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1644511149
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1644511149
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_281
timestamp 1644511149
transform 1 0 26956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1644511149
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_313
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_319
timestamp 1644511149
transform 1 0 30452 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_323
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_343
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1644511149
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_386
timestamp 1644511149
transform 1 0 36616 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_398
timestamp 1644511149
transform 1 0 37720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_405
timestamp 1644511149
transform 1 0 38364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1644511149
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_26
timestamp 1644511149
transform 1 0 3496 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1644511149
transform 1 0 3864 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1644511149
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1644511149
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_67
timestamp 1644511149
transform 1 0 7268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_78
timestamp 1644511149
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_90
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_98
timestamp 1644511149
transform 1 0 10120 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1644511149
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_124
timestamp 1644511149
transform 1 0 12512 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_134
timestamp 1644511149
transform 1 0 13432 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_146
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_190
timestamp 1644511149
transform 1 0 18584 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_198
timestamp 1644511149
transform 1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_207
timestamp 1644511149
transform 1 0 20148 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1644511149
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_257
timestamp 1644511149
transform 1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1644511149
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_288
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_308
timestamp 1644511149
transform 1 0 29440 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_320
timestamp 1644511149
transform 1 0 30544 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1644511149
transform 1 0 3128 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_76
timestamp 1644511149
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_103
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1644511149
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_182
timestamp 1644511149
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_204
timestamp 1644511149
transform 1 0 19872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1644511149
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_261
timestamp 1644511149
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_268
timestamp 1644511149
transform 1 0 25760 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_287
timestamp 1644511149
transform 1 0 27508 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_291
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_349
timestamp 1644511149
transform 1 0 33212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1644511149
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_410
timestamp 1644511149
transform 1 0 38824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1644511149
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_22
timestamp 1644511149
transform 1 0 3128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1644511149
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1644511149
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_78
timestamp 1644511149
transform 1 0 8280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_85
timestamp 1644511149
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_97
timestamp 1644511149
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1644511149
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_152
timestamp 1644511149
transform 1 0 15088 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1644511149
transform 1 0 17296 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_187
timestamp 1644511149
transform 1 0 18308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_306
timestamp 1644511149
transform 1 0 29256 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_326
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_350
timestamp 1644511149
transform 1 0 33304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_357
timestamp 1644511149
transform 1 0 33948 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_377
timestamp 1644511149
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_414
timestamp 1644511149
transform 1 0 39192 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_426
timestamp 1644511149
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1644511149
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1644511149
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_39
timestamp 1644511149
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_51
timestamp 1644511149
transform 1 0 5796 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_63
timestamp 1644511149
transform 1 0 6900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1644511149
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1644511149
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1644511149
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_129
timestamp 1644511149
transform 1 0 12972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1644511149
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_157
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_169
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_315
timestamp 1644511149
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_326
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_336
timestamp 1644511149
transform 1 0 32016 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_344
timestamp 1644511149
transform 1 0 32752 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_368
timestamp 1644511149
transform 1 0 34960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_380
timestamp 1644511149
transform 1 0 36064 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_392
timestamp 1644511149
transform 1 0 37168 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_21
timestamp 1644511149
transform 1 0 3036 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_44
timestamp 1644511149
transform 1 0 5152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1644511149
transform 1 0 9752 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1644511149
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_129
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_141
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_153
timestamp 1644511149
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_176
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1644511149
transform 1 0 18032 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_204
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_254
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_266
timestamp 1644511149
transform 1 0 25576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1644511149
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_313
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_325
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_343
timestamp 1644511149
transform 1 0 32660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_351
timestamp 1644511149
transform 1 0 33396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_380
timestamp 1644511149
transform 1 0 36064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1644511149
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_20
timestamp 1644511149
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1644511149
transform 1 0 4048 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_44
timestamp 1644511149
transform 1 0 5152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_54
timestamp 1644511149
transform 1 0 6072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_64
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1644511149
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_102
timestamp 1644511149
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_114
timestamp 1644511149
transform 1 0 11592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1644511149
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1644511149
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_151
timestamp 1644511149
transform 1 0 14996 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_159
timestamp 1644511149
transform 1 0 15732 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1644511149
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_240
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_280
timestamp 1644511149
transform 1 0 26864 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_292
timestamp 1644511149
transform 1 0 27968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_296
timestamp 1644511149
transform 1 0 28336 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_343
timestamp 1644511149
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_355
timestamp 1644511149
transform 1 0 33764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_63
timestamp 1644511149
transform 1 0 6900 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_75
timestamp 1644511149
transform 1 0 8004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_83
timestamp 1644511149
transform 1 0 8740 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_100
timestamp 1644511149
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_121
timestamp 1644511149
transform 1 0 12236 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_144
timestamp 1644511149
transform 1 0 14352 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1644511149
transform 1 0 15088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_201
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp 1644511149
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1644511149
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1644511149
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_22
timestamp 1644511149
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_45
timestamp 1644511149
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_57
timestamp 1644511149
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_69
timestamp 1644511149
transform 1 0 7452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 1644511149
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_108
timestamp 1644511149
transform 1 0 11040 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_120
timestamp 1644511149
transform 1 0 12144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_174
timestamp 1644511149
transform 1 0 17112 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1644511149
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1644511149
transform 1 0 21804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1644511149
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_6
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_10
timestamp 1644511149
transform 1 0 2024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_73
timestamp 1644511149
transform 1 0 7820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_85
timestamp 1644511149
transform 1 0 8924 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1644511149
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_209
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1644511149
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_16
timestamp 1644511149
transform 1 0 2576 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_50
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_62
timestamp 1644511149
transform 1 0 6808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_74
timestamp 1644511149
transform 1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1644511149
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_13
timestamp 1644511149
transform 1 0 2300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_20
timestamp 1644511149
transform 1 0 2944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_28
timestamp 1644511149
transform 1 0 3680 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_33
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_46
timestamp 1644511149
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1644511149
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_142
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_154
timestamp 1644511149
transform 1 0 15272 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1644511149
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_38
timestamp 1644511149
transform 1 0 4600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_58
timestamp 1644511149
transform 1 0 6440 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_70
timestamp 1644511149
transform 1 0 7544 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1644511149
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1644511149
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1644511149
transform 1 0 10764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_117
timestamp 1644511149
transform 1 0 11868 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_125
timestamp 1644511149
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1644511149
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_161
timestamp 1644511149
transform 1 0 15916 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_25
timestamp 1644511149
transform 1 0 3404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_32
timestamp 1644511149
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_44
timestamp 1644511149
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_66
timestamp 1644511149
transform 1 0 7176 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_74
timestamp 1644511149
transform 1 0 7912 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_101
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_198
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_210
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1644511149
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1644511149
transform 1 0 4048 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1644511149
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_67
timestamp 1644511149
transform 1 0 7268 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1644511149
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_114
timestamp 1644511149
transform 1 0 11592 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_126
timestamp 1644511149
transform 1 0 12696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1644511149
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_170
timestamp 1644511149
transform 1 0 16744 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_182
timestamp 1644511149
transform 1 0 17848 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_7
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_31
timestamp 1644511149
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_43
timestamp 1644511149
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_175
timestamp 1644511149
transform 1 0 17204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_190
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_202
timestamp 1644511149
transform 1 0 19688 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_214
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1644511149
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_64
timestamp 1644511149
transform 1 0 6992 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_76
timestamp 1644511149
transform 1 0 8096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_117
timestamp 1644511149
transform 1 0 11868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_126
timestamp 1644511149
transform 1 0 12696 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1644511149
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_147
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1644511149
transform 1 0 15272 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1644511149
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_174
timestamp 1644511149
transform 1 0 17112 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_19
timestamp 1644511149
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_31
timestamp 1644511149
transform 1 0 3956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_43
timestamp 1644511149
transform 1 0 5060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1644511149
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_73
timestamp 1644511149
transform 1 0 7820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_85
timestamp 1644511149
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_97
timestamp 1644511149
transform 1 0 10028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1644511149
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_129
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_157
timestamp 1644511149
transform 1 0 15548 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 1644511149
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1644511149
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp 1644511149
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_46
timestamp 1644511149
transform 1 0 5336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_54
timestamp 1644511149
transform 1 0 6072 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_63
timestamp 1644511149
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1644511149
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_6
timestamp 1644511149
transform 1 0 1656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_26
timestamp 1644511149
transform 1 0 3496 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1644511149
transform 1 0 4232 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1644511149
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1644511149
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_37
timestamp 1644511149
transform 1 0 4508 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1644511149
transform 1 0 4968 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1644511149
transform 1 0 6072 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1644511149
transform 1 0 7176 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1644511149
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_18
timestamp 1644511149
transform 1 0 2760 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1644511149
transform 1 0 3864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1644511149
transform 1 0 4968 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_14
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_26
timestamp 1644511149
transform 1 0 3496 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_19
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_43
timestamp 1644511149
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_9
timestamp 1644511149
transform 1 0 1932 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_16
timestamp 1644511149
transform 1 0 2576 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_28
timestamp 1644511149
transform 1 0 3680 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_40
timestamp 1644511149
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1644511149
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_14
timestamp 1644511149
transform 1 0 2392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_26
timestamp 1644511149
transform 1 0 3496 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_38
timestamp 1644511149
transform 1 0 4600 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_50
timestamp 1644511149
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_11
timestamp 1644511149
transform 1 0 2116 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_23
timestamp 1644511149
transform 1 0 3220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_31
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_43
timestamp 1644511149
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_7
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_19
timestamp 1644511149
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_340
timestamp 1644511149
transform 1 0 32384 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_352
timestamp 1644511149
transform 1 0 33488 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_364
timestamp 1644511149
transform 1 0 34592 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_376
timestamp 1644511149
transform 1 0 35696 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1644511149
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_33
timestamp 1644511149
transform 1 0 4140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_45
timestamp 1644511149
transform 1 0 5244 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_57
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_69
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1644511149
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_125
timestamp 1644511149
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1644511149
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1644511149
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_200
timestamp 1644511149
transform 1 0 19504 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_212
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1644511149
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_285
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_297
timestamp 1644511149
transform 1 0 28428 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1644511149
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_349
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_353
timestamp 1644511149
transform 1 0 33580 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1644511149
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_393
timestamp 1644511149
transform 1 0 37260 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_405
timestamp 1644511149
transform 1 0 38364 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_417
timestamp 1644511149
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_439
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_447
timestamp 1644511149
transform 1 0 42228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_449
timestamp 1644511149
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_461
timestamp 1644511149
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1644511149
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_505
timestamp 1644511149
transform 1 0 47564 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_517
timestamp 1644511149
transform 1 0 48668 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_561
timestamp 1644511149
transform 1 0 52716 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_573
timestamp 1644511149
transform 1 0 53820 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1644511149
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_597
timestamp 1644511149
transform 1 0 56028 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_603
timestamp 1644511149
transform 1 0 56580 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_615
timestamp 1644511149
transform 1 0 57684 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1644511149
transform 1 0 57868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 53360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1644511149
transform -1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1644511149
transform -1 0 15180 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1644511149
transform 1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4
timestamp 1644511149
transform -1 0 27784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5
timestamp 1644511149
transform 1 0 22816 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_6
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_7
timestamp 1644511149
transform 1 0 32752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_8
timestamp 1644511149
transform -1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_9
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_10
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_11
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_12
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_13
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_14
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_15
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 42320 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 47472 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 52624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0681_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0682_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0683_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0684_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0685_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0686_
timestamp 1644511149
transform 1 0 7360 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0687_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0688_
timestamp 1644511149
transform 1 0 39744 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0689_
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0690_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33212 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0691_
timestamp 1644511149
transform 1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0692_
timestamp 1644511149
transform 1 0 14260 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0693_
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0694_
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0695_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1644511149
transform 1 0 10580 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0700_
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0702_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 1644511149
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _0704_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0705_
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1644511149
transform 1 0 14904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0707_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0708_
timestamp 1644511149
transform 1 0 6440 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0709_
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0710_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_4  _0711_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or3b_1  _0712_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6808 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0713_
timestamp 1644511149
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1644511149
transform 1 0 48484 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0716_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 49312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0717_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0718_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32200 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0719_
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 52164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0721_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 51428 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0722_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50692 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0723_
timestamp 1644511149
transform 1 0 51428 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform 1 0 47564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0725_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50232 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0726_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _0727_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6992 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0728_
timestamp 1644511149
transform 1 0 5520 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0729_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6992 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0730_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0731_
timestamp 1644511149
transform 1 0 6900 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0732_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7820 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0733_
timestamp 1644511149
transform 1 0 6624 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0734_
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0735_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0736_
timestamp 1644511149
transform 1 0 8096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0737_
timestamp 1644511149
transform 1 0 8280 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_4  _0738_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _0739_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33580 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0740_
timestamp 1644511149
transform 1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0741_
timestamp 1644511149
transform 1 0 35972 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0742_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45448 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0744_
timestamp 1644511149
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0745_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0746_
timestamp 1644511149
transform 1 0 29808 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0747_
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0748_
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0749_
timestamp 1644511149
transform 1 0 49864 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_4  _0750_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_4  _0751_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0752_
timestamp 1644511149
transform 1 0 33488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0753_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48852 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0754_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48116 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 1644511149
transform 1 0 47564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1644511149
transform 1 0 50600 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0757_
timestamp 1644511149
transform 1 0 48116 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0758_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 48760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0759_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 49128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0760_
timestamp 1644511149
transform 1 0 50232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0761_
timestamp 1644511149
transform 1 0 47840 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0762_
timestamp 1644511149
transform 1 0 50232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1644511149
transform 1 0 50508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1644511149
transform 1 0 53544 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0765_
timestamp 1644511149
transform 1 0 54372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1644511149
transform 1 0 53636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0767_
timestamp 1644511149
transform 1 0 54648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0768_
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0769_
timestamp 1644511149
transform 1 0 27140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0770_
timestamp 1644511149
transform 1 0 27140 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0771_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 53636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0772_
timestamp 1644511149
transform 1 0 53544 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0773_
timestamp 1644511149
transform 1 0 53728 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0774_
timestamp 1644511149
transform 1 0 55200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0776_
timestamp 1644511149
transform 1 0 51336 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0777_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0778_
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0779_
timestamp 1644511149
transform 1 0 53360 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0780_
timestamp 1644511149
transform 1 0 53636 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0781_
timestamp 1644511149
transform 1 0 54280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0782_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52900 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1644511149
transform 1 0 52992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0784_
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0785_
timestamp 1644511149
transform 1 0 40204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0786_
timestamp 1644511149
transform 1 0 34868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0787_
timestamp 1644511149
transform 1 0 24932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0788_
timestamp 1644511149
transform 1 0 35696 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1644511149
transform 1 0 34408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0790_
timestamp 1644511149
transform 1 0 13248 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0791_
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0792_
timestamp 1644511149
transform 1 0 15272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1644511149
transform 1 0 15088 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0794_
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0795_
timestamp 1644511149
transform 1 0 14996 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0796_
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0797_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0798_
timestamp 1644511149
transform 1 0 11960 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0799_
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _0800_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0801_
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0802_
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0803_
timestamp 1644511149
transform 1 0 21252 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0804_
timestamp 1644511149
transform 1 0 20976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0805_
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0806_
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0807_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0808_
timestamp 1644511149
transform 1 0 13064 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 1644511149
transform 1 0 16652 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0810_
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0811_
timestamp 1644511149
transform 1 0 15732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 1644511149
transform 1 0 21160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0813_
timestamp 1644511149
transform 1 0 20056 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0814_
timestamp 1644511149
transform 1 0 27968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0815_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 1644511149
transform 1 0 19136 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0818_
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0819_
timestamp 1644511149
transform 1 0 13432 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0820_
timestamp 1644511149
transform 1 0 17940 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0821_
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0822_
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0823_
timestamp 1644511149
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0824_
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0825_
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0826_
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0827_
timestamp 1644511149
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0828_
timestamp 1644511149
transform 1 0 15916 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0829_
timestamp 1644511149
transform 1 0 14904 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _0830_
timestamp 1644511149
transform 1 0 12880 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0831_
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0833_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0834_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0835_
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0836_
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0837_
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0838_
timestamp 1644511149
transform 1 0 25760 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0839_
timestamp 1644511149
transform 1 0 12788 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0840_
timestamp 1644511149
transform 1 0 22080 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0841_
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0842_
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0843_
timestamp 1644511149
transform 1 0 16192 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0844_
timestamp 1644511149
transform 1 0 14996 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0845_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0846_
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _0847_
timestamp 1644511149
transform 1 0 35052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0848_
timestamp 1644511149
transform 1 0 25208 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0849_
timestamp 1644511149
transform 1 0 13064 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0851_
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0852_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0853_
timestamp 1644511149
transform 1 0 38548 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0854_
timestamp 1644511149
transform 1 0 37444 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0855_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0856_
timestamp 1644511149
transform 1 0 34040 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0857_
timestamp 1644511149
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0858_
timestamp 1644511149
transform 1 0 46828 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0859_
timestamp 1644511149
transform 1 0 39100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0860_
timestamp 1644511149
transform 1 0 37904 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0861_
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1644511149
transform 1 0 32292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0863_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46368 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _0864_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36156 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0865_
timestamp 1644511149
transform 1 0 36064 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0866_
timestamp 1644511149
transform 1 0 35696 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0867_
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0868_
timestamp 1644511149
transform 1 0 35788 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0869_
timestamp 1644511149
transform 1 0 40020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1644511149
transform 1 0 45080 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1644511149
transform 1 0 46184 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0872_
timestamp 1644511149
transform 1 0 46828 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0873_
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0874_
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0875_
timestamp 1644511149
transform 1 0 36248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0876_
timestamp 1644511149
transform 1 0 40204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0877_
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0878_
timestamp 1644511149
transform 1 0 45356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0879_
timestamp 1644511149
transform 1 0 46460 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0880_
timestamp 1644511149
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0881_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1644511149
transform 1 0 6808 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1644511149
transform 1 0 8648 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0885_
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0886_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7268 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0888_
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0889_
timestamp 1644511149
transform 1 0 35512 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0890_
timestamp 1644511149
transform 1 0 36064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0891_
timestamp 1644511149
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0892_
timestamp 1644511149
transform 1 0 48668 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0893_
timestamp 1644511149
transform 1 0 48760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0895_
timestamp 1644511149
transform 1 0 46920 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0896_
timestamp 1644511149
transform 1 0 45448 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0898_
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0899_
timestamp 1644511149
transform 1 0 45448 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1644511149
transform 1 0 48760 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 1644511149
transform 1 0 48852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0902_
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0903_
timestamp 1644511149
transform 1 0 32108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0904_
timestamp 1644511149
transform 1 0 35052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0905_
timestamp 1644511149
transform 1 0 33488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1644511149
transform 1 0 38548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0907_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0908_
timestamp 1644511149
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0909_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 1644511149
transform 1 0 42320 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1644511149
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0912_
timestamp 1644511149
transform 1 0 41308 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1644511149
transform 1 0 40940 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1644511149
transform 1 0 41308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0915_
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1644511149
transform 1 0 38272 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0918_
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0919_
timestamp 1644511149
transform 1 0 38456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0920_
timestamp 1644511149
transform 1 0 39192 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0921_
timestamp 1644511149
transform 1 0 40756 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1644511149
transform 1 0 40848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0923_
timestamp 1644511149
transform 1 0 41216 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0924_
timestamp 1644511149
transform 1 0 42228 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0925_
timestamp 1644511149
transform 1 0 41124 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0926_
timestamp 1644511149
transform 1 0 31464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0927_
timestamp 1644511149
transform 1 0 35236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0928_
timestamp 1644511149
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0930_
timestamp 1644511149
transform 1 0 40940 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1644511149
transform 1 0 41952 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0932_
timestamp 1644511149
transform 1 0 42688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0933_
timestamp 1644511149
transform 1 0 42228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0934_
timestamp 1644511149
transform 1 0 39928 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1644511149
transform 1 0 41768 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0936_
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0937_
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0938_
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0939_
timestamp 1644511149
transform 1 0 38548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0940_
timestamp 1644511149
transform 1 0 37904 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1644511149
transform 1 0 38916 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1644511149
transform 1 0 38364 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0943_
timestamp 1644511149
transform 1 0 31832 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0944_
timestamp 1644511149
transform 1 0 32108 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1644511149
transform 1 0 31188 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1644511149
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1644511149
transform 1 0 30912 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0948_
timestamp 1644511149
transform 1 0 31004 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0949_
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0950_
timestamp 1644511149
transform 1 0 31096 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 1644511149
transform 1 0 30084 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1644511149
transform 1 0 30176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1644511149
transform 1 0 29532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _0955_
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1644511149
transform 1 0 33028 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0957_
timestamp 1644511149
transform 1 0 33120 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0958_
timestamp 1644511149
transform 1 0 34132 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0960_
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0961_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33856 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0962_
timestamp 1644511149
transform 1 0 33304 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0963_
timestamp 1644511149
transform 1 0 34960 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0964_
timestamp 1644511149
transform 1 0 35696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0965_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35236 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0966_
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0967_
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0968_
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0969_
timestamp 1644511149
transform 1 0 31924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0970_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0973_
timestamp 1644511149
transform 1 0 37076 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0974_
timestamp 1644511149
transform 1 0 20700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1644511149
transform 1 0 26036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0976_
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0977_
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0980_
timestamp 1644511149
transform 1 0 24656 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0981_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0982_
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0984_
timestamp 1644511149
transform 1 0 25576 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0985_
timestamp 1644511149
transform 1 0 44160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0986_
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0987_
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _0988_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32936 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0989_
timestamp 1644511149
transform 1 0 40940 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0990_
timestamp 1644511149
transform 1 0 40572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0992_
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0993_
timestamp 1644511149
transform 1 0 40756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0994_
timestamp 1644511149
transform 1 0 37628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _0995_
timestamp 1644511149
transform 1 0 36984 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0996_
timestamp 1644511149
transform 1 0 40020 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0997_
timestamp 1644511149
transform 1 0 43240 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1644511149
transform 1 0 43516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0999_
timestamp 1644511149
transform 1 0 46828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1000_
timestamp 1644511149
transform 1 0 44068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1001_
timestamp 1644511149
transform 1 0 43240 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1003_
timestamp 1644511149
transform 1 0 36432 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1004_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1005_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 41124 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1006_
timestamp 1644511149
transform 1 0 40756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1008_
timestamp 1644511149
transform 1 0 36064 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1009_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1010_
timestamp 1644511149
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1011_
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1012_
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1013_
timestamp 1644511149
transform 1 0 35144 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _1014_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43792 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1015_
timestamp 1644511149
transform 1 0 44712 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1644511149
transform 1 0 45356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1017_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43792 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp 1644511149
transform 1 0 46184 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1644511149
transform 1 0 46184 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1021_
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1022_
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1023_
timestamp 1644511149
transform 1 0 46184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1024_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 46552 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1644511149
transform 1 0 47932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1026_
timestamp 1644511149
transform 1 0 44528 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1644511149
transform 1 0 43884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1028_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1644511149
transform 1 0 45264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1030_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 43608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1031_
timestamp 1644511149
transform 1 0 41768 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1032_
timestamp 1644511149
transform 1 0 40204 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1034_
timestamp 1644511149
transform 1 0 43516 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1035_
timestamp 1644511149
transform 1 0 42688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1644511149
transform 1 0 42872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1037_
timestamp 1644511149
transform 1 0 33028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1038_
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1039_
timestamp 1644511149
transform 1 0 28612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1040_
timestamp 1644511149
transform 1 0 27416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1041_
timestamp 1644511149
transform 1 0 26680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1042_
timestamp 1644511149
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1043_
timestamp 1644511149
transform 1 0 27600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1044_
timestamp 1644511149
transform 1 0 22448 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1045_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1046_
timestamp 1644511149
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1047_
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1048_
timestamp 1644511149
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1050_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1051_
timestamp 1644511149
transform 1 0 20148 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1052_
timestamp 1644511149
transform 1 0 19964 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1053_
timestamp 1644511149
transform 1 0 19688 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1644511149
transform 1 0 19320 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1644511149
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _1056_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 1644511149
transform 1 0 22080 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1058_
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1059_
timestamp 1644511149
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1060_
timestamp 1644511149
transform 1 0 25300 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1061_
timestamp 1644511149
transform 1 0 25852 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1062_
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1063_
timestamp 1644511149
transform 1 0 20976 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1064_
timestamp 1644511149
transform 1 0 21896 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1065_
timestamp 1644511149
transform 1 0 22724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1066_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1067_
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1644511149
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1069_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1071_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1644511149
transform 1 0 27140 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1073_
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1074_
timestamp 1644511149
transform 1 0 30452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1075_
timestamp 1644511149
transform 1 0 31556 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1077_
timestamp 1644511149
transform 1 0 30544 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1644511149
transform 1 0 31096 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1079_
timestamp 1644511149
transform 1 0 30728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1080_
timestamp 1644511149
transform 1 0 29900 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1083_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1084_
timestamp 1644511149
transform 1 0 32292 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1085_
timestamp 1644511149
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1644511149
transform 1 0 33764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1087_
timestamp 1644511149
transform 1 0 33120 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1088_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1089_
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1644511149
transform 1 0 30544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1093_
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1094_
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1095_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1096_
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1097_
timestamp 1644511149
transform 1 0 31004 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1098_
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1099_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1100_
timestamp 1644511149
transform 1 0 28612 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1101_
timestamp 1644511149
transform 1 0 27140 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1103_
timestamp 1644511149
transform 1 0 30176 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1105_
timestamp 1644511149
transform 1 0 28336 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1106_
timestamp 1644511149
transform 1 0 27600 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1108_
timestamp 1644511149
transform 1 0 32200 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1109_
timestamp 1644511149
transform 1 0 31280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1110_
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1111_
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1112_
timestamp 1644511149
transform 1 0 32660 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1115_
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1644511149
transform 1 0 38732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1644511149
transform 1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1119_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1121_
timestamp 1644511149
transform 1 0 36708 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1122_
timestamp 1644511149
transform 1 0 38732 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1123_
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1124_
timestamp 1644511149
transform 1 0 38732 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1125_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38548 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1126_
timestamp 1644511149
transform 1 0 38272 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1127_
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1128_
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1129_
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1130_
timestamp 1644511149
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1131_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1132_
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1133_
timestamp 1644511149
transform 1 0 13248 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1134_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1135_
timestamp 1644511149
transform 1 0 25392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1136_
timestamp 1644511149
transform 1 0 6900 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1137_
timestamp 1644511149
transform 1 0 7820 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _1138_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_2  _1139_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1140_
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1141_
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1142_
timestamp 1644511149
transform 1 0 17020 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1143_
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand4b_1  _1145_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1644511149
transform 1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1147_
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1148_
timestamp 1644511149
transform 1 0 14444 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1149_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1150_
timestamp 1644511149
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _1151_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8096 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1152_
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1153_
timestamp 1644511149
transform 1 0 14812 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1154_
timestamp 1644511149
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1155_
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _1156_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1157_
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1158_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1159_
timestamp 1644511149
transform 1 0 10580 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1160_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1162_
timestamp 1644511149
transform 1 0 11684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1163_
timestamp 1644511149
transform 1 0 11776 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1164_
timestamp 1644511149
transform 1 0 11408 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1165_
timestamp 1644511149
transform 1 0 9936 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1166_
timestamp 1644511149
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1169_
timestamp 1644511149
transform 1 0 16192 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_2  _1170_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1172_
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1173_
timestamp 1644511149
transform 1 0 12880 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1174_
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1175_
timestamp 1644511149
transform 1 0 17204 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1176_
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1178_
timestamp 1644511149
transform 1 0 12972 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1179_
timestamp 1644511149
transform 1 0 6532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1180_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1181_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1182_
timestamp 1644511149
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1183_
timestamp 1644511149
transform 1 0 14168 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1184_
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1185_
timestamp 1644511149
transform 1 0 16100 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1186_
timestamp 1644511149
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1187_
timestamp 1644511149
transform 1 0 17480 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1188_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1189_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1190_
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1191_
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1192_
timestamp 1644511149
transform 1 0 15548 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1193_
timestamp 1644511149
transform 1 0 6992 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1194_
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1195_
timestamp 1644511149
transform 1 0 17940 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1196_
timestamp 1644511149
transform 1 0 17572 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1197_
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1198_
timestamp 1644511149
transform 1 0 8096 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1199_
timestamp 1644511149
transform 1 0 17848 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1200_
timestamp 1644511149
transform 1 0 28520 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1201_
timestamp 1644511149
transform 1 0 28060 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1202_
timestamp 1644511149
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1203_
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1204_
timestamp 1644511149
transform 1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1205_
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1206_
timestamp 1644511149
transform 1 0 5152 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1207_
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1208_
timestamp 1644511149
transform 1 0 12052 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1209_
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1210_
timestamp 1644511149
transform 1 0 25300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1211_
timestamp 1644511149
transform 1 0 14260 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1212_
timestamp 1644511149
transform 1 0 13248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1213_
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1214_
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1215_
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1216_
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1217_
timestamp 1644511149
transform 1 0 25944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1218_
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1219_
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1220_
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1221_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1222_
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1223_
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1224_
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1225_
timestamp 1644511149
transform 1 0 6624 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1226_
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1227_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1228_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1229_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1230_
timestamp 1644511149
transform 1 0 12420 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1231_
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1232_
timestamp 1644511149
transform 1 0 33580 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1233_
timestamp 1644511149
transform 1 0 32016 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1234_
timestamp 1644511149
transform 1 0 30912 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1235_
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1236_
timestamp 1644511149
transform 1 0 18952 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1237_
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1238_
timestamp 1644511149
transform 1 0 13800 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1239_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1240_
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1644511149
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1242_
timestamp 1644511149
transform 1 0 16836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1243_
timestamp 1644511149
transform 1 0 12420 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1244_
timestamp 1644511149
transform 1 0 32016 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1245_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1246_
timestamp 1644511149
transform 1 0 19504 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1247_
timestamp 1644511149
transform 1 0 19412 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1248_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1249_
timestamp 1644511149
transform 1 0 30912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1250_
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1251_
timestamp 1644511149
transform 1 0 20516 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1252_
timestamp 1644511149
transform 1 0 19044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _1253_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1254_
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1255_
timestamp 1644511149
transform 1 0 33396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1256_
timestamp 1644511149
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1257_
timestamp 1644511149
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1258_
timestamp 1644511149
transform 1 0 19688 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1259_
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1260_
timestamp 1644511149
transform 1 0 18216 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1261_
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1262_
timestamp 1644511149
transform 1 0 15272 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1264_
timestamp 1644511149
transform 1 0 34868 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1265_
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1266_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1267_
timestamp 1644511149
transform 1 0 19320 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1268_
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1269_
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1270_
timestamp 1644511149
transform 1 0 35052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1271_
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1272_
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1273_
timestamp 1644511149
transform 1 0 18124 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1274_
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1275_
timestamp 1644511149
transform 1 0 36156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1276_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1277_
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1278_
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1279_
timestamp 1644511149
transform 1 0 12144 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1280_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35696 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1281_
timestamp 1644511149
transform 1 0 15640 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1282_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1283_
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1284_
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1285_
timestamp 1644511149
transform 1 0 17664 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1286_
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1287_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1288_
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _1289_
timestamp 1644511149
transform 1 0 35972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1290_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1291_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1292_
timestamp 1644511149
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1293_
timestamp 1644511149
transform 1 0 37168 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1294_
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1295_
timestamp 1644511149
transform 1 0 15088 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1296_
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1297_
timestamp 1644511149
transform 1 0 12512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1298_
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1299_
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1300_
timestamp 1644511149
transform 1 0 9752 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1301_
timestamp 1644511149
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1302_
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1303_
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1304_
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1305_
timestamp 1644511149
transform 1 0 15456 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1306_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1307_
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1644511149
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1309_
timestamp 1644511149
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1311_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1644511149
transform 1 0 8832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1313_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _1314_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1315_
timestamp 1644511149
transform 1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1316_
timestamp 1644511149
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1318_
timestamp 1644511149
transform 1 0 2208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1644511149
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1320_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1322_
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1324_
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1326_
timestamp 1644511149
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1327_
timestamp 1644511149
transform 1 0 2760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1328_
timestamp 1644511149
transform 1 0 2852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1329_
timestamp 1644511149
transform 1 0 2208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1330_
timestamp 1644511149
transform 1 0 2668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1331_
timestamp 1644511149
transform 1 0 2392 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1332_
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1333_
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1334_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1335_
timestamp 1644511149
transform 1 0 3312 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1336_
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1337_
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1338_
timestamp 1644511149
transform 1 0 2116 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1339_
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1340_
timestamp 1644511149
transform 1 0 3864 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1341_
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1342_
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1644511149
transform 1 0 2668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1344_
timestamp 1644511149
transform 1 0 2300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1345_
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1346_
timestamp 1644511149
transform 1 0 5060 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1347_
timestamp 1644511149
transform 1 0 5428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1644511149
transform 1 0 3772 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1349_
timestamp 1644511149
transform 1 0 4508 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1644511149
transform 1 0 2300 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1352_
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1353_
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1354_
timestamp 1644511149
transform 1 0 2576 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1355_
timestamp 1644511149
transform 1 0 2300 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1356_
timestamp 1644511149
transform 1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1357_
timestamp 1644511149
transform 1 0 4508 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1358_
timestamp 1644511149
transform 1 0 4692 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1359_
timestamp 1644511149
transform 1 0 6256 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1360_
timestamp 1644511149
transform 1 0 6164 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1361_
timestamp 1644511149
transform 1 0 5612 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1362_
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1644511149
transform 1 0 5152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1364_
timestamp 1644511149
transform 1 0 45080 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1365_
timestamp 1644511149
transform 1 0 52992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1366_
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1367_
timestamp 1644511149
transform 1 0 7912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1368_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1369_
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 1644511149
transform 1 0 10488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1372_
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1373_
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1374_
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1375_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45632 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1376_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 49312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 48760 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 53176 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform 1 0 55844 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 55844 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform 1 0 52992 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 52624 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 14444 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1644511149
transform 1 0 14260 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1644511149
transform 1 0 12880 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform 1 0 15456 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1644511149
transform 1 0 17296 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 21620 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 25392 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1644511149
transform 1 0 21896 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1644511149
transform 1 0 14352 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1644511149
transform 1 0 21528 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1644511149
transform 1 0 46552 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1644511149
transform 1 0 48760 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1644511149
transform 1 0 49128 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1644511149
transform 1 0 50784 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1644511149
transform 1 0 45632 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1644511149
transform 1 0 43976 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1644511149
transform 1 0 41952 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1644511149
transform 1 0 38180 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1644511149
transform 1 0 42964 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1644511149
transform 1 0 43700 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1644511149
transform 1 0 45448 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1644511149
transform 1 0 37904 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1644511149
transform 1 0 29992 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1644511149
transform 1 0 29072 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1644511149
transform 1 0 28244 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1644511149
transform 1 0 31004 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1644511149
transform 1 0 33856 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1434_
timestamp 1644511149
transform 1 0 35236 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1435_
timestamp 1644511149
transform 1 0 35236 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1436_
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1437_
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1438_
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1439_
timestamp 1644511149
transform 1 0 24840 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1440_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1441_
timestamp 1644511149
transform 1 0 26220 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1442_
timestamp 1644511149
transform 1 0 31096 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1443_
timestamp 1644511149
transform 1 0 34500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1444_
timestamp 1644511149
transform 1 0 37352 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1445_
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1446_
timestamp 1644511149
transform 1 0 41124 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1447_
timestamp 1644511149
transform 1 0 28152 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1448_
timestamp 1644511149
transform 1 0 9384 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1449_
timestamp 1644511149
transform 1 0 34776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1450_
timestamp 1644511149
transform 1 0 45264 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1451_
timestamp 1644511149
transform 1 0 46552 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1452_
timestamp 1644511149
transform 1 0 48300 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1453_
timestamp 1644511149
transform 1 0 45448 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1454_
timestamp 1644511149
transform 1 0 40296 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1455_
timestamp 1644511149
transform 1 0 42596 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1456_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1457_
timestamp 1644511149
transform 1 0 23736 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1458_
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1459_
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1460_
timestamp 1644511149
transform 1 0 19596 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1461_
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1462_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1463_
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1464_
timestamp 1644511149
transform 1 0 27232 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1465_
timestamp 1644511149
transform 1 0 30176 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1466_
timestamp 1644511149
transform 1 0 29256 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1467_
timestamp 1644511149
transform 1 0 34132 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1468_
timestamp 1644511149
transform 1 0 31188 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1469_
timestamp 1644511149
transform 1 0 27048 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1470_
timestamp 1644511149
transform 1 0 27968 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1471_
timestamp 1644511149
transform 1 0 28428 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1472_
timestamp 1644511149
transform 1 0 31188 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1473_
timestamp 1644511149
transform 1 0 34592 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1474_
timestamp 1644511149
transform 1 0 37536 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1475_
timestamp 1644511149
transform 1 0 39100 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1476_
timestamp 1644511149
transform 1 0 37904 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1477_
timestamp 1644511149
transform 1 0 40480 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1478_
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1479_
timestamp 1644511149
transform 1 0 10120 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1480_
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1481_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1482_
timestamp 1644511149
transform 1 0 1840 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1483_
timestamp 1644511149
transform 1 0 2576 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1484_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1485_
timestamp 1644511149
transform 1 0 4784 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1486_
timestamp 1644511149
transform 1 0 4232 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1487_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1488_
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1489_
timestamp 1644511149
transform 1 0 4784 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1490_
timestamp 1644511149
transform 1 0 8280 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1491_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1492_
timestamp 1644511149
transform 1 0 10580 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1493_
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1494_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1495_
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1496_
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1497_
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1500_
timestamp 1644511149
transform 1 0 15272 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1501_
timestamp 1644511149
transform 1 0 8188 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1502_
timestamp 1644511149
transform 1 0 10120 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1503_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1504_
timestamp 1644511149
transform 1 0 10764 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1505_
timestamp 1644511149
transform 1 0 8832 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1506_
timestamp 1644511149
transform 1 0 12788 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1507_
timestamp 1644511149
transform 1 0 15548 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1508_
timestamp 1644511149
transform 1 0 16100 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1509_
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1510_
timestamp 1644511149
transform 1 0 13340 0 -1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1511_
timestamp 1644511149
transform 1 0 9108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1512_
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1513_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1514_
timestamp 1644511149
transform 1 0 2024 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1515_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1516_
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1517_
timestamp 1644511149
transform 1 0 2576 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1518_
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1519_
timestamp 1644511149
transform 1 0 1932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1520_
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1521_
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1522_
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1523_
timestamp 1644511149
transform 1 0 1656 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1524_
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1525_
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1526_
timestamp 1644511149
transform 1 0 2116 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1527_
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1528_
timestamp 1644511149
transform 1 0 4968 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1529_
timestamp 1644511149
transform 1 0 1932 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1530_
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1531_
timestamp 1644511149
transform 1 0 2024 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1532_
timestamp 1644511149
transform 1 0 4416 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1533_
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1534_
timestamp 1644511149
transform 1 0 5796 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1535_
timestamp 1644511149
transform 1 0 53360 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1536_
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1537_
timestamp 1644511149
transform 1 0 6072 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1538_
timestamp 1644511149
transform 1 0 9568 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1539_
timestamp 1644511149
transform 1 0 10856 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1540_
timestamp 1644511149
transform 1 0 10396 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1541__183 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1542__184
timestamp 1644511149
transform 1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1543__185
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1544__186
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1545__187
timestamp 1644511149
transform 1 0 13892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1546__179
timestamp 1644511149
transform 1 0 41216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1547__180
timestamp 1644511149
transform 1 0 48760 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1548__181
timestamp 1644511149
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1549__182
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 33672 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 34868 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1644511149
transform 1 0 46460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1644511149
transform 1 0 47932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input18
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input19
timestamp 1644511149
transform 1 0 51060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input20
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input21
timestamp 1644511149
transform 1 0 53912 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input22
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input23
timestamp 1644511149
transform 1 0 56764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input25
timestamp 1644511149
transform 1 0 57684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1644511149
transform 1 0 56856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 2668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 3772 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 2852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  input56 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1472 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 2852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input64
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input65
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input69
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input70 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input72
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 2760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input75
timestamp 1644511149
transform 1 0 1656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1644511149
transform 1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1644511149
transform 1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1644511149
transform 1 0 1472 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1644511149
transform 1 0 3128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1644511149
transform 1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 56212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 35972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 40480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 40388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 45172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1644511149
transform 1 0 49036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1644511149
transform 1 0 50968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1644511149
transform 1 0 51704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1644511149
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1644511149
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1644511149
transform 1 0 55844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1644511149
transform 1 0 23736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1644511149
transform 1 0 2116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1644511149
transform 1 0 2852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1644511149
transform 1 0 2668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1644511149
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3698 41200 3754 42000 6 flash_csb
port 0 nsew signal tristate
rlabel metal2 s 11150 41200 11206 42000 6 flash_io0_read
port 1 nsew signal input
rlabel metal2 s 18694 41200 18750 42000 6 flash_io0_we
port 2 nsew signal tristate
rlabel metal2 s 26146 41200 26202 42000 6 flash_io0_write
port 3 nsew signal tristate
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 4 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 5 nsew signal tristate
rlabel metal2 s 48686 41200 48742 42000 6 flash_io1_write
port 6 nsew signal tristate
rlabel metal2 s 56138 41200 56194 42000 6 flash_sck
port 7 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 8 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 9 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 10 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 11 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 12 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 13 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 14 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 15 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 16 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 17 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 18 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 19 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 20 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 21 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 22 nsew signal tristate
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 23 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 24 nsew signal tristate
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 25 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 26 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 27 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 28 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 29 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 30 nsew signal tristate
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 31 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 32 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 33 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 34 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 35 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 36 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 37 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 38 nsew signal tristate
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 39 nsew signal tristate
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 40 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 41 nsew signal tristate
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 42 nsew signal tristate
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 43 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 44 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 45 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 46 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 47 nsew signal tristate
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 48 nsew signal tristate
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 49 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 50 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 51 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 52 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 53 nsew signal tristate
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 54 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 55 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 56 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 57 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 58 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 59 nsew signal tristate
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 60 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 61 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 62 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 63 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 64 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 65 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 66 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 67 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 68 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 69 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 70 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 71 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 72 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 73 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 74 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 75 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 76 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 77 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 78 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 79 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 80 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 81 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 82 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 83 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 84 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 85 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 86 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 87 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 88 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 89 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 90 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 91 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 92 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 93 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 94 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 95 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 96 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 97 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 98 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 99 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 100 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 101 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 102 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 103 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 104 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 105 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 106 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 107 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 108 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 109 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 110 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 111 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 112 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 113 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 114 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 115 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 116 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 117 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 118 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 119 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 120 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 121 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 122 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 123 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 124 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 125 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 126 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 127 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 128 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 129 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 130 nsew signal tristate
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 131 nsew power input
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 132 nsew ground input
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 132 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 133 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[0]
port 134 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wb_adr_i[10]
port 135 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 136 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 137 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 138 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 139 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[15]
port 140 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[16]
port 141 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[17]
port 142 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_adr_i[18]
port 143 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_adr_i[19]
port 144 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_adr_i[1]
port 145 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_adr_i[20]
port 146 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_adr_i[21]
port 147 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_adr_i[22]
port 148 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[23]
port 149 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_adr_i[2]
port 150 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_adr_i[3]
port 151 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_adr_i[4]
port 152 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 wb_adr_i[5]
port 153 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_adr_i[6]
port 154 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wb_adr_i[7]
port 155 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wb_adr_i[8]
port 156 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wb_adr_i[9]
port 157 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_clk_i
port 158 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wb_cyc_i
port 159 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_data_i[0]
port 160 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_data_i[10]
port 161 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 162 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 163 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 164 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 165 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[15]
port 166 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[16]
port 167 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wb_data_i[17]
port 168 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wb_data_i[18]
port 169 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[19]
port 170 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_data_i[1]
port 171 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[20]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wb_data_i[21]
port 173 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wb_data_i[22]
port 174 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_data_i[23]
port 175 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wb_data_i[24]
port 176 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 wb_data_i[25]
port 177 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[26]
port 178 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wb_data_i[27]
port 179 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_data_i[28]
port 180 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wb_data_i[29]
port 181 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_data_i[2]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 wb_data_i[30]
port 183 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 wb_data_i[31]
port 184 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_data_i[3]
port 185 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_data_i[4]
port 186 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_data_i[5]
port 187 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_data_i[6]
port 188 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_data_i[7]
port 189 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_data_i[8]
port 190 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_data_i[9]
port 191 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_data_o[0]
port 192 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 wb_data_o[10]
port 193 nsew signal tristate
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 194 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 195 nsew signal tristate
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 196 nsew signal tristate
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[14]
port 197 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[15]
port 198 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[16]
port 199 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[17]
port 200 nsew signal tristate
rlabel metal3 s 0 28704 800 28824 6 wb_data_o[18]
port 201 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 wb_data_o[19]
port 202 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 wb_data_o[1]
port 203 nsew signal tristate
rlabel metal3 s 0 31152 800 31272 6 wb_data_o[20]
port 204 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[21]
port 205 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wb_data_o[22]
port 206 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[23]
port 207 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[24]
port 208 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wb_data_o[25]
port 209 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wb_data_o[26]
port 210 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wb_data_o[27]
port 211 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[28]
port 212 nsew signal tristate
rlabel metal3 s 0 39992 800 40112 6 wb_data_o[29]
port 213 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 wb_data_o[2]
port 214 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wb_data_o[30]
port 215 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wb_data_o[31]
port 216 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 wb_data_o[3]
port 217 nsew signal tristate
rlabel metal3 s 0 11024 800 11144 6 wb_data_o[4]
port 218 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 wb_data_o[5]
port 219 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 wb_data_o[6]
port 220 nsew signal tristate
rlabel metal3 s 0 14832 800 14952 6 wb_data_o[7]
port 221 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 wb_data_o[8]
port 222 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 wb_data_o[9]
port 223 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wb_error_o
port 224 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 wb_rst_i
port 225 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wb_sel_i[0]
port 226 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_sel_i[1]
port 227 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_sel_i[2]
port 228 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_sel_i[3]
port 229 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_stall_o
port 230 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 wb_stb_i
port 231 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
<< end >>
