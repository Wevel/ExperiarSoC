magic
tech sky130A
magscale 1 2
timestamp 1653382885
<< viali >>
rect 1593 39593 1627 39627
rect 2329 39593 2363 39627
rect 3985 39593 4019 39627
rect 26433 39593 26467 39627
rect 41429 39593 41463 39627
rect 48973 39593 49007 39627
rect 56425 39593 56459 39627
rect 19257 39457 19291 39491
rect 1409 39389 1443 39423
rect 2145 39389 2179 39423
rect 2881 39389 2915 39423
rect 3065 39253 3099 39287
rect 1409 38913 1443 38947
rect 1593 38709 1627 38743
rect 1593 38505 1627 38539
rect 1409 38301 1443 38335
rect 1409 37825 1443 37859
rect 1593 37621 1627 37655
rect 1409 36737 1443 36771
rect 1593 36601 1627 36635
rect 1409 36125 1443 36159
rect 1593 35989 1627 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 1409 34697 1443 34731
rect 1593 34561 1627 34595
rect 1409 33949 1443 33983
rect 1593 33813 1627 33847
rect 1593 33473 1627 33507
rect 2421 33473 2455 33507
rect 1409 33337 1443 33371
rect 2237 33269 2271 33303
rect 3249 32997 3283 33031
rect 4997 32929 5031 32963
rect 5089 32929 5123 32963
rect 1869 32861 1903 32895
rect 2136 32861 2170 32895
rect 4537 32725 4571 32759
rect 4905 32725 4939 32759
rect 1593 32521 1627 32555
rect 2421 32521 2455 32555
rect 2881 32521 2915 32555
rect 5825 32521 5859 32555
rect 2789 32453 2823 32487
rect 1409 32385 1443 32419
rect 4712 32385 4746 32419
rect 3065 32317 3099 32351
rect 4445 32317 4479 32351
rect 4813 31977 4847 32011
rect 1409 31909 1443 31943
rect 1593 31773 1627 31807
rect 3065 31773 3099 31807
rect 4997 31773 5031 31807
rect 2881 31637 2915 31671
rect 3126 31365 3160 31399
rect 4721 31365 4755 31399
rect 1409 31297 1443 31331
rect 4905 31297 4939 31331
rect 4997 31297 5031 31331
rect 2881 31229 2915 31263
rect 1593 31161 1627 31195
rect 5181 31161 5215 31195
rect 4261 31093 4295 31127
rect 4721 31093 4755 31127
rect 2513 30889 2547 30923
rect 2973 30753 3007 30787
rect 3157 30753 3191 30787
rect 1593 30685 1627 30719
rect 2881 30685 2915 30719
rect 1409 30549 1443 30583
rect 4537 30345 4571 30379
rect 1409 30209 1443 30243
rect 2697 30209 2731 30243
rect 3413 30209 3447 30243
rect 3157 30141 3191 30175
rect 2513 30073 2547 30107
rect 1593 30005 1627 30039
rect 3801 29801 3835 29835
rect 4445 29665 4479 29699
rect 1593 29597 1627 29631
rect 4169 29597 4203 29631
rect 4261 29529 4295 29563
rect 1409 29461 1443 29495
rect 2881 29257 2915 29291
rect 1409 29121 1443 29155
rect 2789 29121 2823 29155
rect 2973 29053 3007 29087
rect 1593 28985 1627 29019
rect 2421 28917 2455 28951
rect 1869 28509 1903 28543
rect 2136 28441 2170 28475
rect 3249 28373 3283 28407
rect 2329 28169 2363 28203
rect 1593 28033 1627 28067
rect 2513 28033 2547 28067
rect 3893 28033 3927 28067
rect 3985 27965 4019 27999
rect 4077 27965 4111 27999
rect 1409 27829 1443 27863
rect 3525 27829 3559 27863
rect 2881 27625 2915 27659
rect 1409 27421 1443 27455
rect 2421 27421 2455 27455
rect 3065 27421 3099 27455
rect 4169 27421 4203 27455
rect 4414 27353 4448 27387
rect 1593 27285 1627 27319
rect 2237 27285 2271 27319
rect 5549 27285 5583 27319
rect 3985 27081 4019 27115
rect 2044 27013 2078 27047
rect 1777 26945 1811 26979
rect 4169 26945 4203 26979
rect 3157 26741 3191 26775
rect 2237 26537 2271 26571
rect 3801 26537 3835 26571
rect 4261 26469 4295 26503
rect 2697 26401 2731 26435
rect 2881 26401 2915 26435
rect 3893 26401 3927 26435
rect 1409 26333 1443 26367
rect 4077 26333 4111 26367
rect 2605 26265 2639 26299
rect 3801 26265 3835 26299
rect 1593 26197 1627 26231
rect 1593 25857 1627 25891
rect 3893 25857 3927 25891
rect 1409 25653 1443 25687
rect 3709 25653 3743 25687
rect 5181 25449 5215 25483
rect 1409 25245 1443 25279
rect 3801 25245 3835 25279
rect 4068 25177 4102 25211
rect 1593 25109 1627 25143
rect 3433 24905 3467 24939
rect 3801 24837 3835 24871
rect 1593 24769 1627 24803
rect 2421 24769 2455 24803
rect 3893 24769 3927 24803
rect 3985 24701 4019 24735
rect 1409 24633 1443 24667
rect 2237 24565 2271 24599
rect 1869 24157 1903 24191
rect 2136 24157 2170 24191
rect 3249 24021 3283 24055
rect 1593 23817 1627 23851
rect 2237 23817 2271 23851
rect 2697 23817 2731 23851
rect 1409 23681 1443 23715
rect 2605 23681 2639 23715
rect 3525 23681 3559 23715
rect 2789 23613 2823 23647
rect 3709 23613 3743 23647
rect 1593 23069 1627 23103
rect 4537 23069 4571 23103
rect 4782 23001 4816 23035
rect 1409 22933 1443 22967
rect 5917 22933 5951 22967
rect 3893 22729 3927 22763
rect 4629 22729 4663 22763
rect 3801 22661 3835 22695
rect 1409 22593 1443 22627
rect 2421 22593 2455 22627
rect 4813 22593 4847 22627
rect 3985 22525 4019 22559
rect 3433 22457 3467 22491
rect 1593 22389 1627 22423
rect 2237 22389 2271 22423
rect 4537 22185 4571 22219
rect 4445 22049 4479 22083
rect 1869 21981 1903 22015
rect 2136 21981 2170 22015
rect 4537 21981 4571 22015
rect 7021 21981 7055 22015
rect 4261 21913 4295 21947
rect 7288 21913 7322 21947
rect 3249 21845 3283 21879
rect 4721 21845 4755 21879
rect 8401 21845 8435 21879
rect 2237 21641 2271 21675
rect 3985 21641 4019 21675
rect 1409 21505 1443 21539
rect 2605 21505 2639 21539
rect 3525 21505 3559 21539
rect 3709 21505 3743 21539
rect 3801 21505 3835 21539
rect 9597 21505 9631 21539
rect 9864 21505 9898 21539
rect 2697 21437 2731 21471
rect 2789 21437 2823 21471
rect 1593 21301 1627 21335
rect 3525 21301 3559 21335
rect 10977 21301 11011 21335
rect 1409 21097 1443 21131
rect 7573 21097 7607 21131
rect 8217 21097 8251 21131
rect 9413 21097 9447 21131
rect 10425 21097 10459 21131
rect 13093 21097 13127 21131
rect 15761 21097 15795 21131
rect 4261 20961 4295 20995
rect 6193 20961 6227 20995
rect 8125 20961 8159 20995
rect 9505 20961 9539 20995
rect 1593 20893 1627 20927
rect 2421 20893 2455 20927
rect 4537 20893 4571 20927
rect 8033 20893 8067 20927
rect 9413 20893 9447 20927
rect 10609 20893 10643 20927
rect 10885 20893 10919 20927
rect 11713 20893 11747 20927
rect 14381 20893 14415 20927
rect 6460 20825 6494 20859
rect 11980 20825 12014 20859
rect 14648 20825 14682 20859
rect 2237 20757 2271 20791
rect 8401 20757 8435 20791
rect 9781 20757 9815 20791
rect 10793 20757 10827 20791
rect 3341 20553 3375 20587
rect 7113 20553 7147 20587
rect 8033 20553 8067 20587
rect 8401 20553 8435 20587
rect 12449 20553 12483 20587
rect 14657 20553 14691 20587
rect 2228 20485 2262 20519
rect 1961 20417 1995 20451
rect 7297 20417 7331 20451
rect 7481 20417 7515 20451
rect 7573 20417 7607 20451
rect 8217 20417 8251 20451
rect 8493 20417 8527 20451
rect 12633 20417 12667 20451
rect 12817 20417 12851 20451
rect 12909 20417 12943 20451
rect 14841 20417 14875 20451
rect 15025 20417 15059 20451
rect 15117 20417 15151 20451
rect 2237 20009 2271 20043
rect 7665 20009 7699 20043
rect 7849 20009 7883 20043
rect 12541 20009 12575 20043
rect 12725 20009 12759 20043
rect 14657 20009 14691 20043
rect 15025 20009 15059 20043
rect 1593 19941 1627 19975
rect 2789 19873 2823 19907
rect 7573 19873 7607 19907
rect 1409 19805 1443 19839
rect 7481 19805 7515 19839
rect 12357 19805 12391 19839
rect 12541 19805 12575 19839
rect 14657 19805 14691 19839
rect 14841 19805 14875 19839
rect 2605 19737 2639 19771
rect 2697 19669 2731 19703
rect 1409 19465 1443 19499
rect 5365 19465 5399 19499
rect 6929 19465 6963 19499
rect 7757 19465 7791 19499
rect 14841 19465 14875 19499
rect 15669 19465 15703 19499
rect 1593 19329 1627 19363
rect 2237 19329 2271 19363
rect 3985 19329 4019 19363
rect 4252 19329 4286 19363
rect 6561 19329 6595 19363
rect 7573 19329 7607 19363
rect 7849 19329 7883 19363
rect 8309 19329 8343 19363
rect 9413 19329 9447 19363
rect 11805 19329 11839 19363
rect 12817 19329 12851 19363
rect 14473 19329 14507 19363
rect 15485 19329 15519 19363
rect 15761 19329 15795 19363
rect 6653 19261 6687 19295
rect 8401 19261 8435 19295
rect 9137 19261 9171 19295
rect 11529 19261 11563 19295
rect 12909 19261 12943 19295
rect 14565 19261 14599 19295
rect 7389 19193 7423 19227
rect 2053 19125 2087 19159
rect 6745 19125 6779 19159
rect 8493 19125 8527 19159
rect 8677 19125 8711 19159
rect 12817 19125 12851 19159
rect 13185 19125 13219 19159
rect 14473 19125 14507 19159
rect 15301 19125 15335 19159
rect 14289 18921 14323 18955
rect 16865 18921 16899 18955
rect 5457 18853 5491 18887
rect 14381 18785 14415 18819
rect 1409 18717 1443 18751
rect 2421 18717 2455 18751
rect 4077 18717 4111 18751
rect 7573 18717 7607 18751
rect 7849 18717 7883 18751
rect 9229 18717 9263 18751
rect 10977 18717 11011 18751
rect 13001 18717 13035 18751
rect 13185 18717 13219 18751
rect 13277 18717 13311 18751
rect 14289 18717 14323 18751
rect 15485 18717 15519 18751
rect 15741 18717 15775 18751
rect 4344 18649 4378 18683
rect 7389 18649 7423 18683
rect 7757 18649 7791 18683
rect 11244 18649 11278 18683
rect 12817 18649 12851 18683
rect 1593 18581 1627 18615
rect 2237 18581 2271 18615
rect 9045 18581 9079 18615
rect 12357 18581 12391 18615
rect 14657 18581 14691 18615
rect 2237 18377 2271 18411
rect 2697 18377 2731 18411
rect 10517 18377 10551 18411
rect 14933 18377 14967 18411
rect 3525 18309 3559 18343
rect 1593 18241 1627 18275
rect 2605 18241 2639 18275
rect 8033 18241 8067 18275
rect 10425 18241 10459 18275
rect 11805 18241 11839 18275
rect 13820 18241 13854 18275
rect 2789 18173 2823 18207
rect 7757 18173 7791 18207
rect 11529 18173 11563 18207
rect 13553 18173 13587 18207
rect 1409 18037 1443 18071
rect 3801 18037 3835 18071
rect 14381 17833 14415 17867
rect 18061 17833 18095 17867
rect 5917 17697 5951 17731
rect 1869 17629 1903 17663
rect 2136 17629 2170 17663
rect 7941 17629 7975 17663
rect 8217 17629 8251 17663
rect 14565 17629 14599 17663
rect 14841 17629 14875 17663
rect 16681 17629 16715 17663
rect 6184 17561 6218 17595
rect 7757 17561 7791 17595
rect 14749 17561 14783 17595
rect 16948 17561 16982 17595
rect 3249 17493 3283 17527
rect 7297 17493 7331 17527
rect 8125 17493 8159 17527
rect 1593 17289 1627 17323
rect 7665 17289 7699 17323
rect 18245 17289 18279 17323
rect 1409 17153 1443 17187
rect 7297 17153 7331 17187
rect 7389 17153 7423 17187
rect 9781 17153 9815 17187
rect 10241 17153 10275 17187
rect 16865 17153 16899 17187
rect 17132 17153 17166 17187
rect 10333 17085 10367 17119
rect 7481 16949 7515 16983
rect 9597 16949 9631 16983
rect 10333 16949 10367 16983
rect 10609 16949 10643 16983
rect 7389 16745 7423 16779
rect 11529 16745 11563 16779
rect 16497 16745 16531 16779
rect 17233 16745 17267 16779
rect 18153 16745 18187 16779
rect 4077 16609 4111 16643
rect 7389 16609 7423 16643
rect 10149 16609 10183 16643
rect 16497 16609 16531 16643
rect 1409 16541 1443 16575
rect 2421 16541 2455 16575
rect 7297 16541 7331 16575
rect 9689 16541 9723 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 12541 16541 12575 16575
rect 16405 16541 16439 16575
rect 17417 16541 17451 16575
rect 17693 16541 17727 16575
rect 18337 16541 18371 16575
rect 18613 16541 18647 16575
rect 4344 16473 4378 16507
rect 10416 16473 10450 16507
rect 12081 16473 12115 16507
rect 18521 16473 18555 16507
rect 1593 16405 1627 16439
rect 2237 16405 2271 16439
rect 5457 16405 5491 16439
rect 7665 16405 7699 16439
rect 9505 16405 9539 16439
rect 16773 16405 16807 16439
rect 17601 16405 17635 16439
rect 7481 16201 7515 16235
rect 7849 16201 7883 16235
rect 17417 16201 17451 16235
rect 2320 16133 2354 16167
rect 1593 16065 1627 16099
rect 2053 16065 2087 16099
rect 6653 16065 6687 16099
rect 6745 16065 6779 16099
rect 7665 16065 7699 16099
rect 7941 16065 7975 16099
rect 10333 16065 10367 16099
rect 10425 16065 10459 16099
rect 11529 16065 11563 16099
rect 11785 16065 11819 16099
rect 13728 16065 13762 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 13461 15997 13495 16031
rect 1409 15861 1443 15895
rect 3433 15861 3467 15895
rect 6837 15861 6871 15895
rect 7021 15861 7055 15895
rect 10333 15861 10367 15895
rect 10701 15861 10735 15895
rect 12909 15861 12943 15895
rect 14841 15861 14875 15895
rect 17049 15861 17083 15895
rect 2145 15657 2179 15691
rect 14473 15657 14507 15691
rect 14841 15657 14875 15691
rect 17233 15657 17267 15691
rect 6653 15589 6687 15623
rect 10793 15589 10827 15623
rect 2605 15521 2639 15555
rect 2697 15521 2731 15555
rect 1593 15453 1627 15487
rect 2513 15453 2547 15487
rect 5273 15453 5307 15487
rect 7665 15453 7699 15487
rect 7849 15453 7883 15487
rect 7941 15453 7975 15487
rect 10977 15453 11011 15487
rect 11161 15453 11195 15487
rect 11253 15453 11287 15487
rect 14473 15453 14507 15487
rect 14657 15453 14691 15487
rect 17233 15453 17267 15487
rect 17417 15453 17451 15487
rect 5540 15385 5574 15419
rect 7481 15385 7515 15419
rect 1409 15317 1443 15351
rect 17601 15317 17635 15351
rect 18613 15113 18647 15147
rect 8309 15045 8343 15079
rect 1409 14977 1443 15011
rect 2421 14977 2455 15011
rect 8125 14977 8159 15011
rect 10057 14977 10091 15011
rect 10241 14977 10275 15011
rect 10333 14977 10367 15011
rect 14197 14977 14231 15011
rect 17500 14977 17534 15011
rect 13921 14909 13955 14943
rect 17233 14909 17267 14943
rect 1593 14841 1627 14875
rect 2237 14773 2271 14807
rect 9873 14773 9907 14807
rect 2329 14569 2363 14603
rect 4353 14569 4387 14603
rect 10333 14569 10367 14603
rect 10885 14569 10919 14603
rect 11253 14569 11287 14603
rect 16681 14569 16715 14603
rect 17509 14569 17543 14603
rect 2789 14433 2823 14467
rect 2973 14433 3007 14467
rect 5825 14433 5859 14467
rect 6009 14433 6043 14467
rect 10977 14433 11011 14467
rect 13553 14433 13587 14467
rect 1593 14365 1627 14399
rect 8953 14365 8987 14399
rect 9220 14365 9254 14399
rect 10885 14365 10919 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 16681 14365 16715 14399
rect 16865 14365 16899 14399
rect 17693 14365 17727 14399
rect 17877 14365 17911 14399
rect 17969 14365 18003 14399
rect 4261 14297 4295 14331
rect 13369 14297 13403 14331
rect 1409 14229 1443 14263
rect 2697 14229 2731 14263
rect 5365 14229 5399 14263
rect 5733 14229 5767 14263
rect 17049 14229 17083 14263
rect 3341 14025 3375 14059
rect 18061 14025 18095 14059
rect 2228 13957 2262 13991
rect 1961 13889 1995 13923
rect 3893 13889 3927 13923
rect 5733 13889 5767 13923
rect 12725 13889 12759 13923
rect 12992 13889 13026 13923
rect 14657 13889 14691 13923
rect 14749 13889 14783 13923
rect 16948 13889 16982 13923
rect 4077 13821 4111 13855
rect 10149 13821 10183 13855
rect 10425 13821 10459 13855
rect 16681 13821 16715 13855
rect 14105 13753 14139 13787
rect 5549 13685 5583 13719
rect 14657 13685 14691 13719
rect 15025 13685 15059 13719
rect 1593 13481 1627 13515
rect 6837 13481 6871 13515
rect 9505 13481 9539 13515
rect 14105 13481 14139 13515
rect 16865 13481 16899 13515
rect 12725 13345 12759 13379
rect 1409 13277 1443 13311
rect 3801 13277 3835 13311
rect 5457 13277 5491 13311
rect 5713 13277 5747 13311
rect 9321 13277 9355 13311
rect 9413 13277 9447 13311
rect 10149 13277 10183 13311
rect 10425 13277 10459 13311
rect 13001 13277 13035 13311
rect 14289 13277 14323 13311
rect 14565 13277 14599 13311
rect 17049 13277 17083 13311
rect 17233 13277 17267 13311
rect 17325 13277 17359 13311
rect 14473 13209 14507 13243
rect 3985 13141 4019 13175
rect 9689 13141 9723 13175
rect 4629 12937 4663 12971
rect 10149 12937 10183 12971
rect 18429 12937 18463 12971
rect 14657 12869 14691 12903
rect 1409 12801 1443 12835
rect 2421 12801 2455 12835
rect 4537 12801 4571 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 8769 12801 8803 12835
rect 9036 12801 9070 12835
rect 10793 12801 10827 12835
rect 13093 12801 13127 12835
rect 14473 12801 14507 12835
rect 15761 12801 15795 12835
rect 15853 12801 15887 12835
rect 17305 12801 17339 12835
rect 4813 12733 4847 12767
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 13369 12733 13403 12767
rect 17049 12733 17083 12767
rect 1593 12597 1627 12631
rect 2237 12597 2271 12631
rect 4169 12597 4203 12631
rect 5641 12597 5675 12631
rect 6377 12597 6411 12631
rect 10885 12597 10919 12631
rect 15761 12597 15795 12631
rect 16129 12597 16163 12631
rect 2237 12393 2271 12427
rect 10149 12393 10183 12427
rect 13093 12393 13127 12427
rect 14289 12393 14323 12427
rect 16957 12393 16991 12427
rect 1409 12325 1443 12359
rect 2789 12257 2823 12291
rect 14197 12257 14231 12291
rect 1593 12189 1627 12223
rect 4537 12189 4571 12223
rect 6285 12189 6319 12223
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 10609 12189 10643 12223
rect 11713 12189 11747 12223
rect 14105 12189 14139 12223
rect 17141 12189 17175 12223
rect 17325 12189 17359 12223
rect 17417 12189 17451 12223
rect 2605 12121 2639 12155
rect 6530 12121 6564 12155
rect 11980 12121 12014 12155
rect 2697 12053 2731 12087
rect 4353 12053 4387 12087
rect 7665 12053 7699 12087
rect 14473 12053 14507 12087
rect 13277 11849 13311 11883
rect 13645 11849 13679 11883
rect 15669 11849 15703 11883
rect 2136 11781 2170 11815
rect 4690 11781 4724 11815
rect 11989 11781 12023 11815
rect 1869 11713 1903 11747
rect 4445 11713 4479 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 13461 11713 13495 11747
rect 13737 11713 13771 11747
rect 15301 11713 15335 11747
rect 16957 11713 16991 11747
rect 15393 11645 15427 11679
rect 17049 11645 17083 11679
rect 3249 11509 3283 11543
rect 5825 11509 5859 11543
rect 8677 11509 8711 11543
rect 12081 11509 12115 11543
rect 15485 11509 15519 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 12817 11305 12851 11339
rect 15945 11305 15979 11339
rect 18705 11305 18739 11339
rect 1593 11237 1627 11271
rect 2145 11237 2179 11271
rect 8953 11169 8987 11203
rect 1409 11101 1443 11135
rect 2329 11101 2363 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 9965 11101 9999 11135
rect 12633 11101 12667 11135
rect 12817 11101 12851 11135
rect 14565 11101 14599 11135
rect 17325 11101 17359 11135
rect 9321 11033 9355 11067
rect 10149 11033 10183 11067
rect 14832 11033 14866 11067
rect 17592 11033 17626 11067
rect 8401 10965 8435 10999
rect 13001 10965 13035 10999
rect 1409 10761 1443 10795
rect 3065 10761 3099 10795
rect 12909 10761 12943 10795
rect 15301 10761 15335 10795
rect 15669 10761 15703 10795
rect 17509 10761 17543 10795
rect 17877 10761 17911 10795
rect 1593 10625 1627 10659
rect 2973 10625 3007 10659
rect 8493 10625 8527 10659
rect 8677 10625 8711 10659
rect 11796 10625 11830 10659
rect 15485 10625 15519 10659
rect 15761 10625 15795 10659
rect 17693 10625 17727 10659
rect 17969 10625 18003 10659
rect 3249 10557 3283 10591
rect 11529 10557 11563 10591
rect 2605 10421 2639 10455
rect 8861 10421 8895 10455
rect 5273 10217 5307 10251
rect 5457 10217 5491 10251
rect 7941 10217 7975 10251
rect 12081 10217 12115 10251
rect 5181 10081 5215 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 2881 10013 2915 10047
rect 4997 10013 5031 10047
rect 5273 10013 5307 10047
rect 6101 10013 6135 10047
rect 8125 10013 8159 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 6368 9945 6402 9979
rect 2697 9877 2731 9911
rect 7481 9877 7515 9911
rect 12449 9877 12483 9911
rect 6377 9673 6411 9707
rect 8953 9673 8987 9707
rect 2780 9605 2814 9639
rect 1409 9537 1443 9571
rect 6561 9537 6595 9571
rect 10057 9537 10091 9571
rect 15761 9537 15795 9571
rect 16937 9537 16971 9571
rect 2513 9469 2547 9503
rect 8493 9469 8527 9503
rect 10333 9469 10367 9503
rect 15853 9469 15887 9503
rect 15945 9469 15979 9503
rect 16681 9469 16715 9503
rect 8861 9401 8895 9435
rect 1593 9333 1627 9367
rect 3893 9333 3927 9367
rect 15393 9333 15427 9367
rect 18061 9333 18095 9367
rect 6009 9129 6043 9163
rect 6193 9129 6227 9163
rect 11989 9129 12023 9163
rect 15945 9129 15979 9163
rect 19257 9129 19291 9163
rect 1409 9061 1443 9095
rect 3249 9061 3283 9095
rect 5641 9061 5675 9095
rect 17693 9061 17727 9095
rect 7573 8993 7607 9027
rect 9137 8993 9171 9027
rect 10057 8993 10091 9027
rect 1593 8925 1627 8959
rect 2237 8925 2271 8959
rect 3065 8925 3099 8959
rect 7849 8925 7883 8959
rect 9229 8925 9263 8959
rect 10609 8925 10643 8959
rect 13369 8925 13403 8959
rect 16129 8925 16163 8959
rect 17877 8925 17911 8959
rect 18153 8925 18187 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 10876 8857 10910 8891
rect 2053 8789 2087 8823
rect 6009 8789 6043 8823
rect 13185 8789 13219 8823
rect 18061 8789 18095 8823
rect 19625 8789 19659 8823
rect 1777 8585 1811 8619
rect 11529 8585 11563 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 17049 8585 17083 8619
rect 19441 8585 19475 8619
rect 2666 8517 2700 8551
rect 6469 8517 6503 8551
rect 7757 8517 7791 8551
rect 8125 8517 8159 8551
rect 13338 8517 13372 8551
rect 19809 8517 19843 8551
rect 20729 8517 20763 8551
rect 1961 8449 1995 8483
rect 2421 8449 2455 8483
rect 6377 8449 6411 8483
rect 7941 8449 7975 8483
rect 10149 8449 10183 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 11989 8449 12023 8483
rect 15853 8449 15887 8483
rect 16129 8449 16163 8483
rect 16681 8449 16715 8483
rect 16865 8449 16899 8483
rect 17141 8449 17175 8483
rect 18153 8449 18187 8483
rect 18429 8449 18463 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 20821 8449 20855 8483
rect 10425 8381 10459 8415
rect 13093 8381 13127 8415
rect 20361 8313 20395 8347
rect 3801 8245 3835 8279
rect 14473 8245 14507 8279
rect 2513 8041 2547 8075
rect 8125 8041 8159 8075
rect 10793 8041 10827 8075
rect 11161 8041 11195 8075
rect 12817 8041 12851 8075
rect 2973 7905 3007 7939
rect 3157 7905 3191 7939
rect 13277 7905 13311 7939
rect 13461 7905 13495 7939
rect 17877 7905 17911 7939
rect 1409 7837 1443 7871
rect 6745 7837 6779 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 17601 7837 17635 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 19717 7837 19751 7871
rect 7012 7769 7046 7803
rect 19257 7769 19291 7803
rect 1593 7701 1627 7735
rect 2881 7701 2915 7735
rect 13185 7701 13219 7735
rect 2145 7497 2179 7531
rect 5181 7497 5215 7531
rect 7113 7497 7147 7531
rect 13461 7497 13495 7531
rect 13829 7497 13863 7531
rect 14933 7497 14967 7531
rect 18797 7497 18831 7531
rect 2605 7429 2639 7463
rect 13093 7429 13127 7463
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 4057 7361 4091 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 8861 7361 8895 7395
rect 10517 7361 10551 7395
rect 10609 7361 10643 7395
rect 12909 7361 12943 7395
rect 13185 7361 13219 7395
rect 13645 7361 13679 7395
rect 13921 7361 13955 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 17417 7361 17451 7395
rect 18613 7361 18647 7395
rect 18889 7361 18923 7395
rect 1961 7293 1995 7327
rect 3801 7293 3835 7327
rect 6653 7293 6687 7327
rect 6745 7293 6779 7327
rect 12725 7293 12759 7327
rect 14565 7293 14599 7327
rect 17141 7293 17175 7327
rect 9229 7225 9263 7259
rect 10517 7157 10551 7191
rect 10885 7157 10919 7191
rect 14289 7157 14323 7191
rect 18429 7157 18463 7191
rect 2881 6953 2915 6987
rect 6101 6953 6135 6987
rect 7389 6953 7423 6987
rect 7297 6885 7331 6919
rect 7205 6817 7239 6851
rect 14289 6817 14323 6851
rect 15853 6817 15887 6851
rect 17141 6817 17175 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 4537 6749 4571 6783
rect 4813 6749 4847 6783
rect 6009 6749 6043 6783
rect 7113 6749 7147 6783
rect 7573 6749 7607 6783
rect 9321 6749 9355 6783
rect 9505 6749 9539 6783
rect 10057 6749 10091 6783
rect 14565 6749 14599 6783
rect 16129 6749 16163 6783
rect 17417 6749 17451 6783
rect 2697 6681 2731 6715
rect 10324 6681 10358 6715
rect 2897 6613 2931 6647
rect 3065 6613 3099 6647
rect 6837 6613 6871 6647
rect 9413 6613 9447 6647
rect 11437 6613 11471 6647
rect 2789 6409 2823 6443
rect 3709 6409 3743 6443
rect 10425 6409 10459 6443
rect 10793 6409 10827 6443
rect 14473 6409 14507 6443
rect 15393 6409 15427 6443
rect 16865 6409 16899 6443
rect 3341 6341 3375 6375
rect 7113 6341 7147 6375
rect 7297 6341 7331 6375
rect 15025 6341 15059 6375
rect 17754 6341 17788 6375
rect 1409 6273 1443 6307
rect 2697 6273 2731 6307
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 15209 6273 15243 6307
rect 15485 6273 15519 6307
rect 17049 6273 17083 6307
rect 14105 6205 14139 6239
rect 17509 6205 17543 6239
rect 1593 6069 1627 6103
rect 18889 6069 18923 6103
rect 14473 5865 14507 5899
rect 15485 5865 15519 5899
rect 16405 5865 16439 5899
rect 3065 5729 3099 5763
rect 6561 5729 6595 5763
rect 16865 5729 16899 5763
rect 16957 5729 16991 5763
rect 1593 5661 1627 5695
rect 3801 5661 3835 5695
rect 6828 5661 6862 5695
rect 14657 5661 14691 5695
rect 14933 5661 14967 5695
rect 15669 5661 15703 5695
rect 15945 5661 15979 5695
rect 2881 5593 2915 5627
rect 14841 5593 14875 5627
rect 1409 5525 1443 5559
rect 2421 5525 2455 5559
rect 2789 5525 2823 5559
rect 7941 5525 7975 5559
rect 15853 5525 15887 5559
rect 16773 5525 16807 5559
rect 1409 5321 1443 5355
rect 3617 5321 3651 5355
rect 4077 5321 4111 5355
rect 12909 5321 12943 5355
rect 14289 5321 14323 5355
rect 15209 5321 15243 5355
rect 16681 5321 16715 5355
rect 18613 5321 18647 5355
rect 14657 5253 14691 5287
rect 15577 5253 15611 5287
rect 17049 5253 17083 5287
rect 18981 5253 19015 5287
rect 1593 5185 1627 5219
rect 2237 5185 2271 5219
rect 2504 5185 2538 5219
rect 4261 5185 4295 5219
rect 4905 5185 4939 5219
rect 6561 5185 6595 5219
rect 9781 5185 9815 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 11785 5185 11819 5219
rect 14473 5185 14507 5219
rect 14749 5185 14783 5219
rect 15393 5185 15427 5219
rect 15669 5185 15703 5219
rect 16865 5185 16899 5219
rect 17141 5185 17175 5219
rect 18797 5185 18831 5219
rect 19073 5185 19107 5219
rect 4721 5117 4755 5151
rect 6377 5117 6411 5151
rect 9873 5117 9907 5151
rect 11529 5117 11563 5151
rect 5089 4981 5123 5015
rect 6745 4981 6779 5015
rect 9965 4981 9999 5015
rect 10149 4981 10183 5015
rect 10609 4981 10643 5015
rect 10977 4981 11011 5015
rect 2421 4777 2455 4811
rect 10333 4777 10367 4811
rect 11161 4777 11195 4811
rect 15393 4777 15427 4811
rect 18245 4777 18279 4811
rect 3801 4641 3835 4675
rect 8953 4641 8987 4675
rect 16589 4641 16623 4675
rect 19257 4641 19291 4675
rect 1409 4573 1443 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4629 4573 4663 4607
rect 5457 4573 5491 4607
rect 6101 4573 6135 4607
rect 6285 4573 6319 4607
rect 11345 4573 11379 4607
rect 11529 4573 11563 4607
rect 11621 4573 11655 4607
rect 15577 4573 15611 4607
rect 15853 4573 15887 4607
rect 16313 4573 16347 4607
rect 18429 4573 18463 4607
rect 18705 4573 18739 4607
rect 19533 4573 19567 4607
rect 24593 4573 24627 4607
rect 9220 4505 9254 4539
rect 15761 4505 15795 4539
rect 1593 4437 1627 4471
rect 3065 4437 3099 4471
rect 4169 4437 4203 4471
rect 6469 4437 6503 4471
rect 18613 4437 18647 4471
rect 24409 4437 24443 4471
rect 10149 4233 10183 4267
rect 6745 4165 6779 4199
rect 18981 4165 19015 4199
rect 19901 4165 19935 4199
rect 1409 4097 1443 4131
rect 2421 4097 2455 4131
rect 3433 4097 3467 4131
rect 3617 4097 3651 4131
rect 3709 4097 3743 4131
rect 4353 4097 4387 4131
rect 5641 4097 5675 4131
rect 6837 4097 6871 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 10241 4097 10275 4131
rect 14289 4097 14323 4131
rect 18613 4097 18647 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19533 4097 19567 4131
rect 19717 4097 19751 4131
rect 19993 4097 20027 4131
rect 6929 4029 6963 4063
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 2237 3961 2271 3995
rect 4997 3961 5031 3995
rect 5457 3961 5491 3995
rect 1593 3893 1627 3927
rect 3249 3893 3283 3927
rect 4169 3893 4203 3927
rect 6377 3893 6411 3927
rect 14105 3893 14139 3927
rect 11253 3689 11287 3723
rect 16589 3689 16623 3723
rect 18245 3689 18279 3723
rect 2605 3621 2639 3655
rect 57989 3621 58023 3655
rect 3801 3553 3835 3587
rect 14657 3553 14691 3587
rect 1685 3485 1719 3519
rect 2421 3485 2455 3519
rect 4057 3485 4091 3519
rect 5825 3485 5859 3519
rect 6469 3485 6503 3519
rect 7113 3485 7147 3519
rect 7757 3485 7791 3519
rect 10701 3485 10735 3519
rect 11437 3485 11471 3519
rect 11621 3485 11655 3519
rect 11713 3485 11747 3519
rect 12633 3485 12667 3519
rect 13553 3485 13587 3519
rect 14933 3485 14967 3519
rect 16129 3485 16163 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 18429 3485 18463 3519
rect 18613 3485 18647 3519
rect 18705 3485 18739 3519
rect 57805 3417 57839 3451
rect 1869 3349 1903 3383
rect 5181 3349 5215 3383
rect 6285 3349 6319 3383
rect 6929 3349 6963 3383
rect 7573 3349 7607 3383
rect 10517 3349 10551 3383
rect 13369 3349 13403 3383
rect 15945 3349 15979 3383
rect 16957 3349 16991 3383
rect 7941 3145 7975 3179
rect 10517 3145 10551 3179
rect 12265 3145 12299 3179
rect 14473 3145 14507 3179
rect 17417 3145 17451 3179
rect 23673 3145 23707 3179
rect 56977 3145 57011 3179
rect 6806 3077 6840 3111
rect 12633 3077 12667 3111
rect 14841 3077 14875 3111
rect 1685 3009 1719 3043
rect 2697 3009 2731 3043
rect 3433 3009 3467 3043
rect 4445 3009 4479 3043
rect 5733 3009 5767 3043
rect 6561 3009 6595 3043
rect 8585 3009 8619 3043
rect 10057 3009 10091 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 12468 3009 12502 3043
rect 12725 3009 12759 3043
rect 13461 3009 13495 3043
rect 14657 3009 14691 3043
rect 14933 3009 14967 3043
rect 16129 3009 16163 3043
rect 17601 3009 17635 3043
rect 17785 3009 17819 3043
rect 17877 3009 17911 3043
rect 19073 3009 19107 3043
rect 19717 3009 19751 3043
rect 21281 3009 21315 3043
rect 23857 3009 23891 3043
rect 33701 3009 33735 3043
rect 56793 3009 56827 3043
rect 1409 2941 1443 2975
rect 4905 2941 4939 2975
rect 13185 2941 13219 2975
rect 33425 2941 33459 2975
rect 4261 2873 4295 2907
rect 9873 2873 9907 2907
rect 15945 2873 15979 2907
rect 19533 2873 19567 2907
rect 21097 2873 21131 2907
rect 2881 2805 2915 2839
rect 3617 2805 3651 2839
rect 5549 2805 5583 2839
rect 8401 2805 8435 2839
rect 9413 2805 9447 2839
rect 11713 2805 11747 2839
rect 16957 2805 16991 2839
rect 18889 2805 18923 2839
rect 20453 2805 20487 2839
rect 22017 2805 22051 2839
rect 25329 2805 25363 2839
rect 32597 2805 32631 2839
rect 35541 2805 35575 2839
rect 37473 2805 37507 2839
rect 39957 2805 39991 2839
rect 42901 2805 42935 2839
rect 44373 2805 44407 2839
rect 47777 2805 47811 2839
rect 50169 2805 50203 2839
rect 53113 2805 53147 2839
rect 54585 2805 54619 2839
rect 58173 2805 58207 2839
rect 10425 2601 10459 2635
rect 25605 2601 25639 2635
rect 27445 2601 27479 2635
rect 28825 2601 28859 2635
rect 30297 2601 30331 2635
rect 32367 2601 32401 2635
rect 45293 2601 45327 2635
rect 16129 2533 16163 2567
rect 21097 2533 21131 2567
rect 54125 2533 54159 2567
rect 2329 2465 2363 2499
rect 5825 2465 5859 2499
rect 14473 2465 14507 2499
rect 16773 2465 16807 2499
rect 1409 2397 1443 2431
rect 3801 2397 3835 2431
rect 5181 2397 5215 2431
rect 6377 2397 6411 2431
rect 8401 2397 8435 2431
rect 9045 2397 9079 2431
rect 10609 2397 10643 2431
rect 10793 2397 10827 2431
rect 10885 2397 10919 2431
rect 11989 2397 12023 2431
rect 13553 2397 13587 2431
rect 14933 2397 14967 2431
rect 16957 2397 16991 2431
rect 17141 2397 17175 2431
rect 17233 2397 17267 2431
rect 17693 2397 17727 2431
rect 18705 2397 18739 2431
rect 19809 2397 19843 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 23121 2397 23155 2431
rect 23857 2397 23891 2431
rect 24685 2397 24719 2431
rect 25789 2397 25823 2431
rect 26433 2397 26467 2431
rect 27629 2397 27663 2431
rect 28273 2397 28307 2431
rect 29009 2397 29043 2431
rect 29745 2397 29779 2431
rect 30481 2397 30515 2431
rect 31125 2397 31159 2431
rect 32137 2397 32171 2431
rect 34069 2397 34103 2431
rect 34897 2397 34931 2431
rect 35173 2397 35207 2431
rect 38117 2397 38151 2431
rect 38761 2397 38795 2431
rect 41889 2397 41923 2431
rect 43085 2397 43119 2431
rect 43637 2397 43671 2431
rect 45109 2397 45143 2431
rect 46029 2397 46063 2431
rect 46581 2397 46615 2431
rect 48053 2397 48087 2431
rect 48973 2397 49007 2431
rect 50169 2397 50203 2431
rect 50997 2397 51031 2431
rect 51917 2397 51951 2431
rect 52745 2397 52779 2431
rect 53941 2397 53975 2431
rect 55321 2397 55355 2431
rect 56241 2397 56275 2431
rect 58081 2397 58115 2431
rect 9781 2329 9815 2363
rect 36461 2329 36495 2363
rect 37933 2329 37967 2363
rect 40325 2329 40359 2363
rect 41044 2329 41078 2363
rect 42901 2329 42935 2363
rect 56977 2329 57011 2363
rect 3985 2261 4019 2295
rect 6561 2261 6595 2295
rect 7573 2261 7607 2295
rect 9229 2261 9263 2295
rect 12173 2261 12207 2295
rect 12725 2261 12759 2295
rect 15117 2261 15151 2295
rect 17877 2261 17911 2295
rect 19993 2261 20027 2295
rect 22385 2261 22419 2295
rect 24869 2261 24903 2295
rect 36553 2261 36587 2295
rect 40417 2261 40451 2295
rect 41153 2261 41187 2295
rect 43821 2261 43855 2295
rect 46765 2261 46799 2295
rect 48237 2261 48271 2295
rect 50353 2261 50387 2295
rect 51181 2261 51215 2295
rect 52929 2261 52963 2295
rect 55505 2261 55539 2295
rect 57069 2261 57103 2295
<< metal1 >>
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1578 39624 1584 39636
rect 1539 39596 1584 39624
rect 1578 39584 1584 39596
rect 1636 39584 1642 39636
rect 2317 39627 2375 39633
rect 2317 39593 2329 39627
rect 2363 39624 2375 39627
rect 2774 39624 2780 39636
rect 2363 39596 2780 39624
rect 2363 39593 2375 39596
rect 2317 39587 2375 39593
rect 2774 39584 2780 39596
rect 2832 39584 2838 39636
rect 3694 39584 3700 39636
rect 3752 39624 3758 39636
rect 3973 39627 4031 39633
rect 3973 39624 3985 39627
rect 3752 39596 3985 39624
rect 3752 39584 3758 39596
rect 3973 39593 3985 39596
rect 4019 39593 4031 39627
rect 3973 39587 4031 39593
rect 26234 39584 26240 39636
rect 26292 39624 26298 39636
rect 26421 39627 26479 39633
rect 26421 39624 26433 39627
rect 26292 39596 26433 39624
rect 26292 39584 26298 39596
rect 26421 39593 26433 39596
rect 26467 39593 26479 39627
rect 41414 39624 41420 39636
rect 41375 39596 41420 39624
rect 26421 39587 26479 39593
rect 41414 39584 41420 39596
rect 41472 39584 41478 39636
rect 48682 39584 48688 39636
rect 48740 39624 48746 39636
rect 48961 39627 49019 39633
rect 48961 39624 48973 39627
rect 48740 39596 48973 39624
rect 48740 39584 48746 39596
rect 48961 39593 48973 39596
rect 49007 39593 49019 39627
rect 48961 39587 49019 39593
rect 56134 39584 56140 39636
rect 56192 39624 56198 39636
rect 56413 39627 56471 39633
rect 56413 39624 56425 39627
rect 56192 39596 56425 39624
rect 56192 39584 56198 39596
rect 56413 39593 56425 39596
rect 56459 39593 56471 39627
rect 56413 39587 56471 39593
rect 18690 39448 18696 39500
rect 18748 39488 18754 39500
rect 19245 39491 19303 39497
rect 19245 39488 19257 39491
rect 18748 39460 19257 39488
rect 18748 39448 18754 39460
rect 19245 39457 19257 39460
rect 19291 39457 19303 39491
rect 19245 39451 19303 39457
rect 1397 39423 1455 39429
rect 1397 39389 1409 39423
rect 1443 39389 1455 39423
rect 2130 39420 2136 39432
rect 2091 39392 2136 39420
rect 1397 39383 1455 39389
rect 1412 39352 1440 39383
rect 2130 39380 2136 39392
rect 2188 39380 2194 39432
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39420 2927 39423
rect 6638 39420 6644 39432
rect 2915 39392 6644 39420
rect 2915 39389 2927 39392
rect 2869 39383 2927 39389
rect 6638 39380 6644 39392
rect 6696 39380 6702 39432
rect 2314 39352 2320 39364
rect 1412 39324 2320 39352
rect 2314 39312 2320 39324
rect 2372 39312 2378 39364
rect 3050 39284 3056 39296
rect 3011 39256 3056 39284
rect 3050 39244 3056 39256
rect 3108 39244 3114 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 2498 38944 2504 38956
rect 1443 38916 2504 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 2498 38904 2504 38916
rect 2556 38904 2562 38956
rect 1578 38740 1584 38752
rect 1539 38712 1584 38740
rect 1578 38700 1584 38712
rect 1636 38700 1642 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1486 38496 1492 38548
rect 1544 38536 1550 38548
rect 1581 38539 1639 38545
rect 1581 38536 1593 38539
rect 1544 38508 1593 38536
rect 1544 38496 1550 38508
rect 1581 38505 1593 38508
rect 1627 38505 1639 38539
rect 1581 38499 1639 38505
rect 1397 38335 1455 38341
rect 1397 38301 1409 38335
rect 1443 38332 1455 38335
rect 1486 38332 1492 38344
rect 1443 38304 1492 38332
rect 1443 38301 1455 38304
rect 1397 38295 1455 38301
rect 1486 38292 1492 38304
rect 1544 38292 1550 38344
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 1670 37856 1676 37868
rect 1443 37828 1676 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1670 37816 1676 37828
rect 1728 37816 1734 37868
rect 1578 37652 1584 37664
rect 1539 37624 1584 37652
rect 1578 37612 1584 37624
rect 1636 37612 1642 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1762 36768 1768 36780
rect 1443 36740 1768 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1762 36728 1768 36740
rect 1820 36728 1826 36780
rect 1578 36632 1584 36644
rect 1539 36604 1584 36632
rect 1578 36592 1584 36604
rect 1636 36592 1642 36644
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36156 1455 36159
rect 1854 36156 1860 36168
rect 1443 36128 1860 36156
rect 1443 36125 1455 36128
rect 1397 36119 1455 36125
rect 1854 36116 1860 36128
rect 1912 36116 1918 36168
rect 1578 36020 1584 36032
rect 1539 35992 1584 36020
rect 1578 35980 1584 35992
rect 1636 35980 1642 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1946 35068 1952 35080
rect 1443 35040 1952 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1946 35028 1952 35040
rect 2004 35028 2010 35080
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1397 34731 1455 34737
rect 1397 34697 1409 34731
rect 1443 34728 1455 34731
rect 2866 34728 2872 34740
rect 1443 34700 2872 34728
rect 1443 34697 1455 34700
rect 1397 34691 1455 34697
rect 2866 34688 2872 34700
rect 2924 34688 2930 34740
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33980 1455 33983
rect 6270 33980 6276 33992
rect 1443 33952 6276 33980
rect 1443 33949 1455 33952
rect 1397 33943 1455 33949
rect 6270 33940 6276 33952
rect 6328 33940 6334 33992
rect 1578 33844 1584 33856
rect 1539 33816 1584 33844
rect 1578 33804 1584 33816
rect 1636 33804 1642 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1578 33504 1584 33516
rect 1539 33476 1584 33504
rect 1578 33464 1584 33476
rect 1636 33464 1642 33516
rect 2406 33504 2412 33516
rect 2367 33476 2412 33504
rect 2406 33464 2412 33476
rect 2464 33464 2470 33516
rect 1397 33371 1455 33377
rect 1397 33337 1409 33371
rect 1443 33368 1455 33371
rect 4982 33368 4988 33380
rect 1443 33340 4988 33368
rect 1443 33337 1455 33340
rect 1397 33331 1455 33337
rect 4982 33328 4988 33340
rect 5040 33328 5046 33380
rect 2130 33260 2136 33312
rect 2188 33300 2194 33312
rect 2225 33303 2283 33309
rect 2225 33300 2237 33303
rect 2188 33272 2237 33300
rect 2188 33260 2194 33272
rect 2225 33269 2237 33272
rect 2271 33269 2283 33303
rect 2225 33263 2283 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 3237 33031 3295 33037
rect 3237 32997 3249 33031
rect 3283 33028 3295 33031
rect 4614 33028 4620 33040
rect 3283 33000 4620 33028
rect 3283 32997 3295 33000
rect 3237 32991 3295 32997
rect 4614 32988 4620 33000
rect 4672 32988 4678 33040
rect 4982 32960 4988 32972
rect 4943 32932 4988 32960
rect 4982 32920 4988 32932
rect 5040 32920 5046 32972
rect 5074 32920 5080 32972
rect 5132 32960 5138 32972
rect 5132 32932 5177 32960
rect 5132 32920 5138 32932
rect 2130 32901 2136 32904
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32861 1915 32895
rect 2124 32892 2136 32901
rect 2091 32864 2136 32892
rect 1857 32855 1915 32861
rect 2124 32855 2136 32864
rect 1872 32824 1900 32855
rect 2130 32852 2136 32855
rect 2188 32852 2194 32904
rect 2774 32824 2780 32836
rect 1872 32796 2780 32824
rect 2774 32784 2780 32796
rect 2832 32784 2838 32836
rect 4525 32759 4583 32765
rect 4525 32725 4537 32759
rect 4571 32756 4583 32759
rect 4798 32756 4804 32768
rect 4571 32728 4804 32756
rect 4571 32725 4583 32728
rect 4525 32719 4583 32725
rect 4798 32716 4804 32728
rect 4856 32716 4862 32768
rect 4890 32716 4896 32768
rect 4948 32756 4954 32768
rect 4948 32728 4993 32756
rect 4948 32716 4954 32728
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1578 32552 1584 32564
rect 1539 32524 1584 32552
rect 1578 32512 1584 32524
rect 1636 32512 1642 32564
rect 2406 32552 2412 32564
rect 2367 32524 2412 32552
rect 2406 32512 2412 32524
rect 2464 32512 2470 32564
rect 2866 32552 2872 32564
rect 2827 32524 2872 32552
rect 2866 32512 2872 32524
rect 2924 32512 2930 32564
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 5813 32555 5871 32561
rect 5813 32552 5825 32555
rect 4948 32524 5825 32552
rect 4948 32512 4954 32524
rect 5813 32521 5825 32524
rect 5859 32521 5871 32555
rect 5813 32515 5871 32521
rect 2777 32487 2835 32493
rect 2777 32453 2789 32487
rect 2823 32484 2835 32487
rect 4614 32484 4620 32496
rect 2823 32456 4620 32484
rect 2823 32453 2835 32456
rect 2777 32447 2835 32453
rect 4614 32444 4620 32456
rect 4672 32444 4678 32496
rect 4706 32425 4712 32428
rect 1397 32419 1455 32425
rect 1397 32385 1409 32419
rect 1443 32385 1455 32419
rect 1397 32379 1455 32385
rect 4700 32379 4712 32425
rect 4764 32416 4770 32428
rect 4764 32388 4800 32416
rect 1412 32212 1440 32379
rect 4706 32376 4712 32379
rect 4764 32376 4770 32388
rect 3053 32351 3111 32357
rect 3053 32317 3065 32351
rect 3099 32348 3111 32351
rect 3142 32348 3148 32360
rect 3099 32320 3148 32348
rect 3099 32317 3111 32320
rect 3053 32311 3111 32317
rect 3142 32308 3148 32320
rect 3200 32308 3206 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 2774 32240 2780 32292
rect 2832 32280 2838 32292
rect 4448 32280 4476 32311
rect 2832 32252 4476 32280
rect 2832 32240 2838 32252
rect 7558 32212 7564 32224
rect 1412 32184 7564 32212
rect 7558 32172 7564 32184
rect 7616 32172 7622 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 4706 31968 4712 32020
rect 4764 32008 4770 32020
rect 4801 32011 4859 32017
rect 4801 32008 4813 32011
rect 4764 31980 4813 32008
rect 4764 31968 4770 31980
rect 4801 31977 4813 31980
rect 4847 31977 4859 32011
rect 4801 31971 4859 31977
rect 1397 31943 1455 31949
rect 1397 31909 1409 31943
rect 1443 31940 1455 31943
rect 2958 31940 2964 31952
rect 1443 31912 2964 31940
rect 1443 31909 1455 31912
rect 1397 31903 1455 31909
rect 2958 31900 2964 31912
rect 3016 31900 3022 31952
rect 1578 31804 1584 31816
rect 1539 31776 1584 31804
rect 1578 31764 1584 31776
rect 1636 31764 1642 31816
rect 3050 31804 3056 31816
rect 3011 31776 3056 31804
rect 3050 31764 3056 31776
rect 3108 31764 3114 31816
rect 4798 31764 4804 31816
rect 4856 31804 4862 31816
rect 4985 31807 5043 31813
rect 4985 31804 4997 31807
rect 4856 31776 4997 31804
rect 4856 31764 4862 31776
rect 4985 31773 4997 31776
rect 5031 31773 5043 31807
rect 4985 31767 5043 31773
rect 2866 31668 2872 31680
rect 2827 31640 2872 31668
rect 2866 31628 2872 31640
rect 2924 31628 2930 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2866 31356 2872 31408
rect 2924 31396 2930 31408
rect 3114 31399 3172 31405
rect 3114 31396 3126 31399
rect 2924 31368 3126 31396
rect 2924 31356 2930 31368
rect 3114 31365 3126 31368
rect 3160 31365 3172 31399
rect 3114 31359 3172 31365
rect 4614 31356 4620 31408
rect 4672 31396 4678 31408
rect 4709 31399 4767 31405
rect 4709 31396 4721 31399
rect 4672 31368 4721 31396
rect 4672 31356 4678 31368
rect 4709 31365 4721 31368
rect 4755 31365 4767 31399
rect 4709 31359 4767 31365
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31328 1455 31331
rect 3418 31328 3424 31340
rect 1443 31300 3424 31328
rect 1443 31297 1455 31300
rect 1397 31291 1455 31297
rect 3418 31288 3424 31300
rect 3476 31288 3482 31340
rect 4890 31328 4896 31340
rect 4851 31300 4896 31328
rect 4890 31288 4896 31300
rect 4948 31288 4954 31340
rect 4982 31288 4988 31340
rect 5040 31328 5046 31340
rect 5040 31300 5085 31328
rect 5040 31288 5046 31300
rect 2774 31220 2780 31272
rect 2832 31260 2838 31272
rect 2869 31263 2927 31269
rect 2869 31260 2881 31263
rect 2832 31232 2881 31260
rect 2832 31220 2838 31232
rect 2869 31229 2881 31232
rect 2915 31229 2927 31263
rect 2869 31223 2927 31229
rect 1578 31192 1584 31204
rect 1539 31164 1584 31192
rect 1578 31152 1584 31164
rect 1636 31152 1642 31204
rect 4614 31152 4620 31204
rect 4672 31192 4678 31204
rect 5169 31195 5227 31201
rect 5169 31192 5181 31195
rect 4672 31164 5181 31192
rect 4672 31152 4678 31164
rect 5169 31161 5181 31164
rect 5215 31161 5227 31195
rect 5169 31155 5227 31161
rect 2866 31084 2872 31136
rect 2924 31124 2930 31136
rect 4249 31127 4307 31133
rect 4249 31124 4261 31127
rect 2924 31096 4261 31124
rect 2924 31084 2930 31096
rect 4249 31093 4261 31096
rect 4295 31124 4307 31127
rect 4709 31127 4767 31133
rect 4709 31124 4721 31127
rect 4295 31096 4721 31124
rect 4295 31093 4307 31096
rect 4249 31087 4307 31093
rect 4709 31093 4721 31096
rect 4755 31093 4767 31127
rect 4709 31087 4767 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 2501 30923 2559 30929
rect 2501 30889 2513 30923
rect 2547 30920 2559 30923
rect 3050 30920 3056 30932
rect 2547 30892 3056 30920
rect 2547 30889 2559 30892
rect 2501 30883 2559 30889
rect 3050 30880 3056 30892
rect 3108 30880 3114 30932
rect 2958 30784 2964 30796
rect 2919 30756 2964 30784
rect 2958 30744 2964 30756
rect 3016 30744 3022 30796
rect 3142 30744 3148 30796
rect 3200 30784 3206 30796
rect 4890 30784 4896 30796
rect 3200 30756 4896 30784
rect 3200 30744 3206 30756
rect 4890 30744 4896 30756
rect 4948 30784 4954 30796
rect 5074 30784 5080 30796
rect 4948 30756 5080 30784
rect 4948 30744 4954 30756
rect 5074 30744 5080 30756
rect 5132 30744 5138 30796
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 2866 30716 2872 30728
rect 2827 30688 2872 30716
rect 2866 30676 2872 30688
rect 2924 30676 2930 30728
rect 1397 30583 1455 30589
rect 1397 30549 1409 30583
rect 1443 30580 1455 30583
rect 4706 30580 4712 30592
rect 1443 30552 4712 30580
rect 1443 30549 1455 30552
rect 1397 30543 1455 30549
rect 4706 30540 4712 30552
rect 4764 30540 4770 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 4525 30379 4583 30385
rect 4525 30345 4537 30379
rect 4571 30376 4583 30379
rect 4982 30376 4988 30388
rect 4571 30348 4988 30376
rect 4571 30345 4583 30348
rect 4525 30339 4583 30345
rect 4982 30336 4988 30348
rect 5040 30336 5046 30388
rect 7742 30308 7748 30320
rect 1412 30280 7748 30308
rect 1412 30249 1440 30280
rect 7742 30268 7748 30280
rect 7800 30268 7806 30320
rect 1397 30243 1455 30249
rect 1397 30209 1409 30243
rect 1443 30209 1455 30243
rect 2682 30240 2688 30252
rect 2643 30212 2688 30240
rect 1397 30203 1455 30209
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 3401 30243 3459 30249
rect 3401 30240 3413 30243
rect 2976 30212 3413 30240
rect 2976 30172 3004 30212
rect 3401 30209 3413 30212
rect 3447 30209 3459 30243
rect 3401 30203 3459 30209
rect 2516 30144 3004 30172
rect 3145 30175 3203 30181
rect 2516 30113 2544 30144
rect 3145 30141 3157 30175
rect 3191 30141 3203 30175
rect 3145 30135 3203 30141
rect 2501 30107 2559 30113
rect 2501 30073 2513 30107
rect 2547 30073 2559 30107
rect 2501 30067 2559 30073
rect 2774 30064 2780 30116
rect 2832 30104 2838 30116
rect 2958 30104 2964 30116
rect 2832 30076 2964 30104
rect 2832 30064 2838 30076
rect 2958 30064 2964 30076
rect 3016 30104 3022 30116
rect 3160 30104 3188 30135
rect 3016 30076 3188 30104
rect 3016 30064 3022 30076
rect 1578 30036 1584 30048
rect 1539 30008 1584 30036
rect 1578 29996 1584 30008
rect 1636 29996 1642 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2682 29792 2688 29844
rect 2740 29832 2746 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 2740 29804 3801 29832
rect 2740 29792 2746 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 4433 29699 4491 29705
rect 4433 29665 4445 29699
rect 4479 29696 4491 29699
rect 4890 29696 4896 29708
rect 4479 29668 4896 29696
rect 4479 29665 4491 29668
rect 4433 29659 4491 29665
rect 4890 29656 4896 29668
rect 4948 29656 4954 29708
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29628 4215 29631
rect 4982 29628 4988 29640
rect 4203 29600 4988 29628
rect 4203 29597 4215 29600
rect 4157 29591 4215 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 4249 29563 4307 29569
rect 4249 29529 4261 29563
rect 4295 29560 4307 29563
rect 4706 29560 4712 29572
rect 4295 29532 4712 29560
rect 4295 29529 4307 29532
rect 4249 29523 4307 29529
rect 4706 29520 4712 29532
rect 4764 29520 4770 29572
rect 1397 29495 1455 29501
rect 1397 29461 1409 29495
rect 1443 29492 1455 29495
rect 2866 29492 2872 29504
rect 1443 29464 2872 29492
rect 1443 29461 1455 29464
rect 1397 29455 1455 29461
rect 2866 29452 2872 29464
rect 2924 29452 2930 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 2866 29288 2872 29300
rect 2827 29260 2872 29288
rect 2866 29248 2872 29260
rect 2924 29248 2930 29300
rect 7650 29220 7656 29232
rect 1412 29192 7656 29220
rect 1412 29161 1440 29192
rect 7650 29180 7656 29192
rect 7708 29180 7714 29232
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29121 1455 29155
rect 2774 29152 2780 29164
rect 2735 29124 2780 29152
rect 1397 29115 1455 29121
rect 2774 29112 2780 29124
rect 2832 29112 2838 29164
rect 2682 29044 2688 29096
rect 2740 29084 2746 29096
rect 2961 29087 3019 29093
rect 2961 29084 2973 29087
rect 2740 29056 2973 29084
rect 2740 29044 2746 29056
rect 2961 29053 2973 29056
rect 3007 29053 3019 29087
rect 2961 29047 3019 29053
rect 1578 29016 1584 29028
rect 1539 28988 1584 29016
rect 1578 28976 1584 28988
rect 1636 28976 1642 29028
rect 2409 28951 2467 28957
rect 2409 28917 2421 28951
rect 2455 28948 2467 28951
rect 2498 28948 2504 28960
rect 2455 28920 2504 28948
rect 2455 28917 2467 28920
rect 2409 28911 2467 28917
rect 2498 28908 2504 28920
rect 2556 28908 2562 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1857 28543 1915 28549
rect 1857 28509 1869 28543
rect 1903 28540 1915 28543
rect 2958 28540 2964 28552
rect 1903 28512 2964 28540
rect 1903 28509 1915 28512
rect 1857 28503 1915 28509
rect 2958 28500 2964 28512
rect 3016 28500 3022 28552
rect 2124 28475 2182 28481
rect 2124 28441 2136 28475
rect 2170 28472 2182 28475
rect 2314 28472 2320 28484
rect 2170 28444 2320 28472
rect 2170 28441 2182 28444
rect 2124 28435 2182 28441
rect 2314 28432 2320 28444
rect 2372 28432 2378 28484
rect 2774 28364 2780 28416
rect 2832 28404 2838 28416
rect 3237 28407 3295 28413
rect 3237 28404 3249 28407
rect 2832 28376 3249 28404
rect 2832 28364 2838 28376
rect 3237 28373 3249 28376
rect 3283 28404 3295 28407
rect 3786 28404 3792 28416
rect 3283 28376 3792 28404
rect 3283 28373 3295 28376
rect 3237 28367 3295 28373
rect 3786 28364 3792 28376
rect 3844 28364 3850 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2314 28200 2320 28212
rect 2275 28172 2320 28200
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 1394 28024 1400 28076
rect 1452 28064 1458 28076
rect 1581 28067 1639 28073
rect 1581 28064 1593 28067
rect 1452 28036 1593 28064
rect 1452 28024 1458 28036
rect 1581 28033 1593 28036
rect 1627 28033 1639 28067
rect 2498 28064 2504 28076
rect 2459 28036 2504 28064
rect 1581 28027 1639 28033
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2590 28024 2596 28076
rect 2648 28024 2654 28076
rect 3878 28064 3884 28076
rect 3839 28036 3884 28064
rect 3878 28024 3884 28036
rect 3936 28024 3942 28076
rect 2498 27888 2504 27940
rect 2556 27928 2562 27940
rect 2608 27928 2636 28024
rect 2682 27956 2688 28008
rect 2740 27956 2746 28008
rect 3970 27996 3976 28008
rect 3931 27968 3976 27996
rect 3970 27956 3976 27968
rect 4028 27956 4034 28008
rect 4065 27999 4123 28005
rect 4065 27965 4077 27999
rect 4111 27965 4123 27999
rect 4065 27959 4123 27965
rect 2556 27900 2636 27928
rect 2700 27928 2728 27956
rect 4080 27928 4108 27959
rect 2700 27900 4108 27928
rect 2556 27888 2562 27900
rect 1397 27863 1455 27869
rect 1397 27829 1409 27863
rect 1443 27860 1455 27863
rect 2682 27860 2688 27872
rect 1443 27832 2688 27860
rect 1443 27829 1455 27832
rect 1397 27823 1455 27829
rect 2682 27820 2688 27832
rect 2740 27820 2746 27872
rect 3513 27863 3571 27869
rect 3513 27829 3525 27863
rect 3559 27860 3571 27863
rect 4062 27860 4068 27872
rect 3559 27832 4068 27860
rect 3559 27829 3571 27832
rect 3513 27823 3571 27829
rect 4062 27820 4068 27832
rect 4120 27820 4126 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 2869 27659 2927 27665
rect 2869 27625 2881 27659
rect 2915 27656 2927 27659
rect 3970 27656 3976 27668
rect 2915 27628 3976 27656
rect 2915 27625 2927 27628
rect 2869 27619 2927 27625
rect 3970 27616 3976 27628
rect 4028 27616 4034 27668
rect 1412 27492 4292 27520
rect 1412 27461 1440 27492
rect 1397 27455 1455 27461
rect 1397 27421 1409 27455
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 2314 27412 2320 27464
rect 2372 27452 2378 27464
rect 2409 27455 2467 27461
rect 2409 27452 2421 27455
rect 2372 27424 2421 27452
rect 2372 27412 2378 27424
rect 2409 27421 2421 27424
rect 2455 27421 2467 27455
rect 3050 27452 3056 27464
rect 3011 27424 3056 27452
rect 2409 27415 2467 27421
rect 3050 27412 3056 27424
rect 3108 27412 3114 27464
rect 3694 27452 3700 27464
rect 3160 27424 3700 27452
rect 2958 27344 2964 27396
rect 3016 27384 3022 27396
rect 3160 27384 3188 27424
rect 3694 27412 3700 27424
rect 3752 27452 3758 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 3752 27424 4169 27452
rect 3752 27412 3758 27424
rect 4157 27421 4169 27424
rect 4203 27421 4215 27455
rect 4264 27452 4292 27492
rect 13078 27452 13084 27464
rect 4264 27424 13084 27452
rect 4157 27415 4215 27421
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 3016 27356 3188 27384
rect 3016 27344 3022 27356
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 4402 27387 4460 27393
rect 4402 27384 4414 27387
rect 4028 27356 4414 27384
rect 4028 27344 4034 27356
rect 4402 27353 4414 27356
rect 4448 27353 4460 27387
rect 4402 27347 4460 27353
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 2222 27316 2228 27328
rect 2183 27288 2228 27316
rect 2222 27276 2228 27288
rect 2280 27276 2286 27328
rect 3878 27276 3884 27328
rect 3936 27316 3942 27328
rect 5537 27319 5595 27325
rect 5537 27316 5549 27319
rect 3936 27288 5549 27316
rect 3936 27276 3942 27288
rect 5537 27285 5549 27288
rect 5583 27285 5595 27319
rect 5537 27279 5595 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 3970 27112 3976 27124
rect 3931 27084 3976 27112
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 2032 27047 2090 27053
rect 2032 27013 2044 27047
rect 2078 27044 2090 27047
rect 2222 27044 2228 27056
rect 2078 27016 2228 27044
rect 2078 27013 2090 27016
rect 2032 27007 2090 27013
rect 2222 27004 2228 27016
rect 2280 27004 2286 27056
rect 1765 26979 1823 26985
rect 1765 26945 1777 26979
rect 1811 26976 1823 26979
rect 2958 26976 2964 26988
rect 1811 26948 2964 26976
rect 1811 26945 1823 26948
rect 1765 26939 1823 26945
rect 2958 26936 2964 26948
rect 3016 26936 3022 26988
rect 4154 26976 4160 26988
rect 4115 26948 4160 26976
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 3142 26772 3148 26784
rect 3103 26744 3148 26772
rect 3142 26732 3148 26744
rect 3200 26732 3206 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 2225 26571 2283 26577
rect 2225 26537 2237 26571
rect 2271 26568 2283 26571
rect 2314 26568 2320 26580
rect 2271 26540 2320 26568
rect 2271 26537 2283 26540
rect 2225 26531 2283 26537
rect 2314 26528 2320 26540
rect 2372 26528 2378 26580
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 3789 26571 3847 26577
rect 3789 26568 3801 26571
rect 3200 26540 3801 26568
rect 3200 26528 3206 26540
rect 3789 26537 3801 26540
rect 3835 26537 3847 26571
rect 3789 26531 3847 26537
rect 4249 26503 4307 26509
rect 1412 26472 4200 26500
rect 1412 26373 1440 26472
rect 2682 26392 2688 26444
rect 2740 26432 2746 26444
rect 2740 26404 2785 26432
rect 2740 26392 2746 26404
rect 2866 26392 2872 26444
rect 2924 26432 2930 26444
rect 3878 26432 3884 26444
rect 2924 26404 2969 26432
rect 3839 26404 3884 26432
rect 2924 26392 2930 26404
rect 3878 26392 3884 26404
rect 3936 26392 3942 26444
rect 4172 26432 4200 26472
rect 4249 26469 4261 26503
rect 4295 26500 4307 26503
rect 4706 26500 4712 26512
rect 4295 26472 4712 26500
rect 4295 26469 4307 26472
rect 4249 26463 4307 26469
rect 4706 26460 4712 26472
rect 4764 26460 4770 26512
rect 15746 26432 15752 26444
rect 4172 26404 15752 26432
rect 15746 26392 15752 26404
rect 15804 26392 15810 26444
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 3970 26324 3976 26376
rect 4028 26364 4034 26376
rect 4065 26367 4123 26373
rect 4065 26364 4077 26367
rect 4028 26336 4077 26364
rect 4028 26324 4034 26336
rect 4065 26333 4077 26336
rect 4111 26333 4123 26367
rect 4065 26327 4123 26333
rect 2593 26299 2651 26305
rect 2593 26265 2605 26299
rect 2639 26296 2651 26299
rect 3142 26296 3148 26308
rect 2639 26268 3148 26296
rect 2639 26265 2651 26268
rect 2593 26259 2651 26265
rect 3142 26256 3148 26268
rect 3200 26256 3206 26308
rect 3786 26296 3792 26308
rect 3747 26268 3792 26296
rect 3786 26256 3792 26268
rect 3844 26256 3850 26308
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 3878 25888 3884 25900
rect 3839 25860 3884 25888
rect 3878 25848 3884 25860
rect 3936 25848 3942 25900
rect 1397 25687 1455 25693
rect 1397 25653 1409 25687
rect 1443 25684 1455 25687
rect 3602 25684 3608 25696
rect 1443 25656 3608 25684
rect 1443 25653 1455 25656
rect 1397 25647 1455 25653
rect 3602 25644 3608 25656
rect 3660 25644 3666 25696
rect 3697 25687 3755 25693
rect 3697 25653 3709 25687
rect 3743 25684 3755 25687
rect 4062 25684 4068 25696
rect 3743 25656 4068 25684
rect 3743 25653 3755 25656
rect 3697 25647 3755 25653
rect 4062 25644 4068 25656
rect 4120 25644 4126 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 5169 25483 5227 25489
rect 5169 25480 5181 25483
rect 4028 25452 5181 25480
rect 4028 25440 4034 25452
rect 5169 25449 5181 25452
rect 5215 25449 5227 25483
rect 5169 25443 5227 25449
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 1412 25208 1440 25239
rect 2774 25236 2780 25288
rect 2832 25276 2838 25288
rect 3694 25276 3700 25288
rect 2832 25248 3700 25276
rect 2832 25236 2838 25248
rect 3694 25236 3700 25248
rect 3752 25276 3758 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3752 25248 3801 25276
rect 3752 25236 3758 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 12250 25276 12256 25288
rect 3789 25239 3847 25245
rect 3988 25248 12256 25276
rect 3988 25208 4016 25248
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 4062 25217 4068 25220
rect 1412 25180 4016 25208
rect 4056 25171 4068 25217
rect 4120 25208 4126 25220
rect 4120 25180 4156 25208
rect 4062 25168 4068 25171
rect 4120 25168 4126 25180
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 3421 24939 3479 24945
rect 3421 24905 3433 24939
rect 3467 24936 3479 24939
rect 3878 24936 3884 24948
rect 3467 24908 3884 24936
rect 3467 24905 3479 24908
rect 3421 24899 3479 24905
rect 3878 24896 3884 24908
rect 3936 24896 3942 24948
rect 3789 24871 3847 24877
rect 3789 24837 3801 24871
rect 3835 24868 3847 24871
rect 3970 24868 3976 24880
rect 3835 24840 3976 24868
rect 3835 24837 3847 24840
rect 3789 24831 3847 24837
rect 3970 24828 3976 24840
rect 4028 24828 4034 24880
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 2222 24760 2228 24812
rect 2280 24800 2286 24812
rect 2409 24803 2467 24809
rect 2409 24800 2421 24803
rect 2280 24772 2421 24800
rect 2280 24760 2286 24772
rect 2409 24769 2421 24772
rect 2455 24769 2467 24803
rect 2409 24763 2467 24769
rect 3602 24760 3608 24812
rect 3660 24800 3666 24812
rect 3881 24803 3939 24809
rect 3881 24800 3893 24803
rect 3660 24772 3893 24800
rect 3660 24760 3666 24772
rect 3881 24769 3893 24772
rect 3927 24769 3939 24803
rect 3881 24763 3939 24769
rect 2590 24692 2596 24744
rect 2648 24732 2654 24744
rect 3973 24735 4031 24741
rect 3973 24732 3985 24735
rect 2648 24704 3985 24732
rect 2648 24692 2654 24704
rect 3973 24701 3985 24704
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 1397 24667 1455 24673
rect 1397 24633 1409 24667
rect 1443 24664 1455 24667
rect 2682 24664 2688 24676
rect 1443 24636 2688 24664
rect 1443 24633 1455 24636
rect 1397 24627 1455 24633
rect 2682 24624 2688 24636
rect 2740 24624 2746 24676
rect 2130 24556 2136 24608
rect 2188 24596 2194 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 2188 24568 2237 24596
rect 2188 24556 2194 24568
rect 2225 24565 2237 24568
rect 2271 24565 2283 24599
rect 2225 24559 2283 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 2130 24197 2136 24200
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 2124 24188 2136 24197
rect 2091 24160 2136 24188
rect 1857 24151 1915 24157
rect 2124 24151 2136 24160
rect 1872 24120 1900 24151
rect 2130 24148 2136 24151
rect 2188 24148 2194 24200
rect 2774 24120 2780 24132
rect 1872 24092 2780 24120
rect 2774 24080 2780 24092
rect 2832 24080 2838 24132
rect 1394 24012 1400 24064
rect 1452 24052 1458 24064
rect 1762 24052 1768 24064
rect 1452 24024 1768 24052
rect 1452 24012 1458 24024
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 1854 24012 1860 24064
rect 1912 24052 1918 24064
rect 2130 24052 2136 24064
rect 1912 24024 2136 24052
rect 1912 24012 1918 24024
rect 2130 24012 2136 24024
rect 2188 24012 2194 24064
rect 3237 24055 3295 24061
rect 3237 24021 3249 24055
rect 3283 24052 3295 24055
rect 3326 24052 3332 24064
rect 3283 24024 3332 24052
rect 3283 24021 3295 24024
rect 3237 24015 3295 24021
rect 3326 24012 3332 24024
rect 3384 24012 3390 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 2222 23848 2228 23860
rect 2183 23820 2228 23848
rect 2222 23808 2228 23820
rect 2280 23808 2286 23860
rect 2682 23848 2688 23860
rect 2643 23820 2688 23848
rect 2682 23808 2688 23820
rect 2740 23808 2746 23860
rect 1397 23715 1455 23721
rect 1397 23681 1409 23715
rect 1443 23712 1455 23715
rect 1854 23712 1860 23724
rect 1443 23684 1860 23712
rect 1443 23681 1455 23684
rect 1397 23675 1455 23681
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23712 2651 23715
rect 3326 23712 3332 23724
rect 2639 23684 3332 23712
rect 2639 23681 2651 23684
rect 2593 23675 2651 23681
rect 3326 23672 3332 23684
rect 3384 23672 3390 23724
rect 3510 23712 3516 23724
rect 3471 23684 3516 23712
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 2682 23604 2688 23656
rect 2740 23644 2746 23656
rect 2777 23647 2835 23653
rect 2777 23644 2789 23647
rect 2740 23616 2789 23644
rect 2740 23604 2746 23616
rect 2777 23613 2789 23616
rect 2823 23644 2835 23647
rect 3697 23647 3755 23653
rect 3697 23644 3709 23647
rect 2823 23616 3709 23644
rect 2823 23613 2835 23616
rect 2777 23607 2835 23613
rect 3697 23613 3709 23616
rect 3743 23613 3755 23647
rect 3697 23607 3755 23613
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 4062 23100 4068 23112
rect 2832 23072 4068 23100
rect 2832 23060 2838 23072
rect 4062 23060 4068 23072
rect 4120 23100 4126 23112
rect 4525 23103 4583 23109
rect 4525 23100 4537 23103
rect 4120 23072 4537 23100
rect 4120 23060 4126 23072
rect 4525 23069 4537 23072
rect 4571 23069 4583 23103
rect 4525 23063 4583 23069
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 4770 23035 4828 23041
rect 4770 23032 4782 23035
rect 4672 23004 4782 23032
rect 4672 22992 4678 23004
rect 4770 23001 4782 23004
rect 4816 23001 4828 23035
rect 4770 22995 4828 23001
rect 1397 22967 1455 22973
rect 1397 22933 1409 22967
rect 1443 22964 1455 22967
rect 3878 22964 3884 22976
rect 1443 22936 3884 22964
rect 1443 22933 1455 22936
rect 1397 22927 1455 22933
rect 3878 22924 3884 22936
rect 3936 22924 3942 22976
rect 3970 22924 3976 22976
rect 4028 22964 4034 22976
rect 5905 22967 5963 22973
rect 5905 22964 5917 22967
rect 4028 22936 5917 22964
rect 4028 22924 4034 22936
rect 5905 22933 5917 22936
rect 5951 22933 5963 22967
rect 5905 22927 5963 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1486 22720 1492 22772
rect 1544 22760 1550 22772
rect 1946 22760 1952 22772
rect 1544 22732 1952 22760
rect 1544 22720 1550 22732
rect 1946 22720 1952 22732
rect 2004 22720 2010 22772
rect 3878 22760 3884 22772
rect 3839 22732 3884 22760
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 4614 22760 4620 22772
rect 4575 22732 4620 22760
rect 4614 22720 4620 22732
rect 4672 22720 4678 22772
rect 3694 22652 3700 22704
rect 3752 22692 3758 22704
rect 3789 22695 3847 22701
rect 3789 22692 3801 22695
rect 3752 22664 3801 22692
rect 3752 22652 3758 22664
rect 3789 22661 3801 22664
rect 3835 22692 3847 22695
rect 3970 22692 3976 22704
rect 3835 22664 3976 22692
rect 3835 22661 3847 22664
rect 3789 22655 3847 22661
rect 3970 22652 3976 22664
rect 4028 22652 4034 22704
rect 1397 22627 1455 22633
rect 1397 22593 1409 22627
rect 1443 22624 1455 22627
rect 1486 22624 1492 22636
rect 1443 22596 1492 22624
rect 1443 22593 1455 22596
rect 1397 22587 1455 22593
rect 1486 22584 1492 22596
rect 1544 22584 1550 22636
rect 2406 22624 2412 22636
rect 2367 22596 2412 22624
rect 2406 22584 2412 22596
rect 2464 22584 2470 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 2590 22516 2596 22568
rect 2648 22556 2654 22568
rect 3973 22559 4031 22565
rect 3973 22556 3985 22559
rect 2648 22528 3985 22556
rect 2648 22516 2654 22528
rect 3973 22525 3985 22528
rect 4019 22525 4031 22559
rect 3973 22519 4031 22525
rect 3421 22491 3479 22497
rect 3421 22457 3433 22491
rect 3467 22488 3479 22491
rect 4816 22488 4844 22587
rect 3467 22460 4844 22488
rect 3467 22457 3479 22460
rect 3421 22451 3479 22457
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 2130 22380 2136 22432
rect 2188 22420 2194 22432
rect 2225 22423 2283 22429
rect 2225 22420 2237 22423
rect 2188 22392 2237 22420
rect 2188 22380 2194 22392
rect 2225 22389 2237 22392
rect 2271 22389 2283 22423
rect 2225 22383 2283 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 4525 22219 4583 22225
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 5442 22216 5448 22228
rect 4571 22188 5448 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 4120 22120 5488 22148
rect 4120 22108 4126 22120
rect 4433 22083 4491 22089
rect 4433 22049 4445 22083
rect 4479 22080 4491 22083
rect 4706 22080 4712 22092
rect 4479 22052 4712 22080
rect 4479 22049 4491 22052
rect 4433 22043 4491 22049
rect 4706 22040 4712 22052
rect 4764 22040 4770 22092
rect 5460 22080 5488 22120
rect 5460 22052 5672 22080
rect 2130 22021 2136 22024
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 21981 1915 22015
rect 2124 22012 2136 22021
rect 2091 21984 2136 22012
rect 1857 21975 1915 21981
rect 2124 21975 2136 21984
rect 1872 21944 1900 21975
rect 2130 21972 2136 21975
rect 2188 21972 2194 22024
rect 3970 21972 3976 22024
rect 4028 22012 4034 22024
rect 4525 22015 4583 22021
rect 4525 22012 4537 22015
rect 4028 21984 4537 22012
rect 4028 21972 4034 21984
rect 4525 21981 4537 21984
rect 4571 21981 4583 22015
rect 5644 22012 5672 22052
rect 6178 22012 6184 22024
rect 5644 21984 6184 22012
rect 4525 21975 4583 21981
rect 6178 21972 6184 21984
rect 6236 22012 6242 22024
rect 7009 22015 7067 22021
rect 7009 22012 7021 22015
rect 6236 21984 7021 22012
rect 6236 21972 6242 21984
rect 7009 21981 7021 21984
rect 7055 22012 7067 22015
rect 9674 22012 9680 22024
rect 7055 21984 9680 22012
rect 7055 21981 7067 21984
rect 7009 21975 7067 21981
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 2774 21944 2780 21956
rect 1872 21916 2780 21944
rect 2774 21904 2780 21916
rect 2832 21904 2838 21956
rect 4249 21947 4307 21953
rect 4249 21913 4261 21947
rect 4295 21944 4307 21947
rect 4798 21944 4804 21956
rect 4295 21916 4804 21944
rect 4295 21913 4307 21916
rect 4249 21907 4307 21913
rect 4798 21904 4804 21916
rect 4856 21904 4862 21956
rect 7276 21947 7334 21953
rect 7276 21913 7288 21947
rect 7322 21944 7334 21947
rect 8018 21944 8024 21956
rect 7322 21916 8024 21944
rect 7322 21913 7334 21916
rect 7276 21907 7334 21913
rect 8018 21904 8024 21916
rect 8076 21904 8082 21956
rect 3234 21876 3240 21888
rect 3195 21848 3240 21876
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 4706 21876 4712 21888
rect 4667 21848 4712 21876
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 8110 21876 8116 21888
rect 6328 21848 8116 21876
rect 6328 21836 6334 21848
rect 8110 21836 8116 21848
rect 8168 21876 8174 21888
rect 8389 21879 8447 21885
rect 8389 21876 8401 21879
rect 8168 21848 8401 21876
rect 8168 21836 8174 21848
rect 8389 21845 8401 21848
rect 8435 21845 8447 21879
rect 8389 21839 8447 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 2406 21672 2412 21684
rect 2271 21644 2412 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 3970 21672 3976 21684
rect 3931 21644 3976 21672
rect 3970 21632 3976 21644
rect 4028 21632 4034 21684
rect 17310 21604 17316 21616
rect 1412 21576 17316 21604
rect 1412 21545 1440 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21536 2651 21539
rect 3234 21536 3240 21548
rect 2639 21508 3240 21536
rect 2639 21505 2651 21508
rect 2593 21499 2651 21505
rect 2682 21468 2688 21480
rect 2643 21440 2688 21468
rect 2682 21428 2688 21440
rect 2740 21428 2746 21480
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21437 2835 21471
rect 2777 21431 2835 21437
rect 2590 21360 2596 21412
rect 2648 21400 2654 21412
rect 2792 21400 2820 21431
rect 2648 21372 2820 21400
rect 2648 21360 2654 21372
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 2884 21332 2912 21508
rect 3234 21496 3240 21508
rect 3292 21496 3298 21548
rect 3326 21496 3332 21548
rect 3384 21536 3390 21548
rect 3513 21539 3571 21545
rect 3513 21536 3525 21539
rect 3384 21508 3525 21536
rect 3384 21496 3390 21508
rect 3513 21505 3525 21508
rect 3559 21505 3571 21539
rect 3694 21536 3700 21548
rect 3655 21508 3700 21536
rect 3513 21499 3571 21505
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 3786 21496 3792 21548
rect 3844 21536 3850 21548
rect 9585 21539 9643 21545
rect 3844 21508 3889 21536
rect 3844 21496 3850 21508
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9674 21536 9680 21548
rect 9631 21508 9680 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9674 21496 9680 21508
rect 9732 21496 9738 21548
rect 9852 21539 9910 21545
rect 9852 21505 9864 21539
rect 9898 21536 9910 21539
rect 10410 21536 10416 21548
rect 9898 21508 10416 21536
rect 9898 21505 9910 21508
rect 9852 21499 9910 21505
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 3513 21335 3571 21341
rect 3513 21332 3525 21335
rect 2884 21304 3525 21332
rect 3513 21301 3525 21304
rect 3559 21301 3571 21335
rect 10962 21332 10968 21344
rect 10923 21304 10968 21332
rect 3513 21295 3571 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1397 21131 1455 21137
rect 1397 21097 1409 21131
rect 1443 21128 1455 21131
rect 2682 21128 2688 21140
rect 1443 21100 2688 21128
rect 1443 21097 1455 21100
rect 1397 21091 1455 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 7558 21128 7564 21140
rect 7519 21100 7564 21128
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 8205 21131 8263 21137
rect 8205 21097 8217 21131
rect 8251 21128 8263 21131
rect 9398 21128 9404 21140
rect 8251 21100 9404 21128
rect 8251 21097 8263 21100
rect 8205 21091 8263 21097
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 10410 21128 10416 21140
rect 10371 21100 10416 21128
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 15746 21128 15752 21140
rect 15707 21100 15752 21128
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 7742 21020 7748 21072
rect 7800 21060 7806 21072
rect 10962 21060 10968 21072
rect 7800 21032 10968 21060
rect 7800 21020 7806 21032
rect 4249 20995 4307 21001
rect 4249 20961 4261 20995
rect 4295 20992 4307 20995
rect 4706 20992 4712 21004
rect 4295 20964 4712 20992
rect 4295 20961 4307 20964
rect 4249 20955 4307 20961
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 6178 20992 6184 21004
rect 6139 20964 6184 20992
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 8110 20992 8116 21004
rect 8071 20964 8116 20992
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 9508 21001 9536 21032
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 9950 20952 9956 21004
rect 10008 20992 10014 21004
rect 10008 20964 10916 20992
rect 10008 20952 10014 20964
rect 1394 20884 1400 20936
rect 1452 20924 1458 20936
rect 1581 20927 1639 20933
rect 1581 20924 1593 20927
rect 1452 20896 1593 20924
rect 1452 20884 1458 20896
rect 1581 20893 1593 20896
rect 1627 20893 1639 20927
rect 2406 20924 2412 20936
rect 2367 20896 2412 20924
rect 1581 20887 1639 20893
rect 2406 20884 2412 20896
rect 2464 20884 2470 20936
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 8021 20927 8079 20933
rect 4571 20896 4752 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 4724 20868 4752 20896
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8294 20924 8300 20936
rect 8067 20896 8300 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 8294 20884 8300 20896
rect 8352 20924 8358 20936
rect 9401 20927 9459 20933
rect 9401 20924 9413 20927
rect 8352 20896 9413 20924
rect 8352 20884 8358 20896
rect 9401 20893 9413 20896
rect 9447 20893 9459 20927
rect 10594 20924 10600 20936
rect 10555 20896 10600 20924
rect 9401 20887 9459 20893
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10888 20933 10916 20964
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20893 10931 20927
rect 10873 20887 10931 20893
rect 10962 20884 10968 20936
rect 11020 20924 11026 20936
rect 11701 20927 11759 20933
rect 11701 20924 11713 20927
rect 11020 20896 11713 20924
rect 11020 20884 11026 20896
rect 11701 20893 11713 20896
rect 11747 20893 11759 20927
rect 12526 20924 12532 20936
rect 11701 20887 11759 20893
rect 11808 20896 12532 20924
rect 4706 20816 4712 20868
rect 4764 20816 4770 20868
rect 6448 20859 6506 20865
rect 6448 20825 6460 20859
rect 6494 20856 6506 20859
rect 7098 20856 7104 20868
rect 6494 20828 7104 20856
rect 6494 20825 6506 20828
rect 6448 20819 6506 20825
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 10612 20856 10640 20884
rect 11808 20856 11836 20896
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 10612 20828 11836 20856
rect 11968 20859 12026 20865
rect 11968 20825 11980 20859
rect 12014 20856 12026 20859
rect 12434 20856 12440 20868
rect 12014 20828 12440 20856
rect 12014 20825 12026 20828
rect 11968 20819 12026 20825
rect 12434 20816 12440 20828
rect 12492 20816 12498 20868
rect 2222 20788 2228 20800
rect 2183 20760 2228 20788
rect 2222 20748 2228 20760
rect 2280 20748 2286 20800
rect 8386 20788 8392 20800
rect 8347 20760 8392 20788
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 9769 20791 9827 20797
rect 9769 20757 9781 20791
rect 9815 20788 9827 20791
rect 10781 20791 10839 20797
rect 10781 20788 10793 20791
rect 9815 20760 10793 20788
rect 9815 20757 9827 20760
rect 9769 20751 9827 20757
rect 10781 20757 10793 20760
rect 10827 20757 10839 20791
rect 10781 20751 10839 20757
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 14384 20788 14412 20887
rect 14642 20865 14648 20868
rect 14636 20819 14648 20865
rect 14700 20856 14706 20868
rect 14700 20828 14736 20856
rect 14642 20816 14648 20819
rect 14700 20816 14706 20828
rect 11020 20760 14412 20788
rect 11020 20748 11026 20760
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 3326 20584 3332 20596
rect 3239 20556 3332 20584
rect 3326 20544 3332 20556
rect 3384 20584 3390 20596
rect 3786 20584 3792 20596
rect 3384 20556 3792 20584
rect 3384 20544 3390 20556
rect 3786 20544 3792 20556
rect 3844 20544 3850 20596
rect 7098 20584 7104 20596
rect 7059 20556 7104 20584
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 7466 20544 7472 20596
rect 7524 20584 7530 20596
rect 8018 20584 8024 20596
rect 7524 20556 7604 20584
rect 7979 20556 8024 20584
rect 7524 20544 7530 20556
rect 2222 20525 2228 20528
rect 2216 20516 2228 20525
rect 2183 20488 2228 20516
rect 2216 20479 2228 20488
rect 2222 20476 2228 20479
rect 2280 20476 2286 20528
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2774 20448 2780 20460
rect 1995 20420 2780 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 7576 20457 7604 20556
rect 8018 20544 8024 20556
rect 8076 20544 8082 20596
rect 8386 20584 8392 20596
rect 8347 20556 8392 20584
rect 8386 20544 8392 20556
rect 8444 20544 8450 20596
rect 12434 20584 12440 20596
rect 12395 20556 12440 20584
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 14642 20584 14648 20596
rect 14603 20556 14648 20584
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 12636 20488 14872 20516
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20448 7343 20451
rect 7469 20451 7527 20457
rect 7331 20420 7420 20448
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 7392 20312 7420 20420
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20448 8539 20451
rect 8570 20448 8576 20460
rect 8527 20420 8576 20448
rect 8527 20417 8539 20420
rect 8481 20411 8539 20417
rect 7484 20380 7512 20411
rect 7834 20380 7840 20392
rect 7484 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 7650 20312 7656 20324
rect 7392 20284 7656 20312
rect 7650 20272 7656 20284
rect 7708 20312 7714 20324
rect 8220 20312 8248 20411
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 12526 20408 12532 20460
rect 12584 20448 12590 20460
rect 12636 20457 12664 20488
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12584 20420 12633 20448
rect 12584 20408 12590 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12768 20420 12817 20448
rect 12768 20408 12774 20420
rect 12805 20417 12817 20420
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 12897 20451 12955 20457
rect 12897 20417 12909 20451
rect 12943 20448 12955 20451
rect 13538 20448 13544 20460
rect 12943 20420 13544 20448
rect 12943 20417 12955 20420
rect 12897 20411 12955 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 14844 20457 14872 20488
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20417 14887 20451
rect 15010 20448 15016 20460
rect 14971 20420 15016 20448
rect 14829 20411 14887 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15160 20420 15205 20448
rect 15160 20408 15166 20420
rect 7708 20284 8248 20312
rect 7708 20272 7714 20284
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 2225 20043 2283 20049
rect 2225 20009 2237 20043
rect 2271 20040 2283 20043
rect 2406 20040 2412 20052
rect 2271 20012 2412 20040
rect 2271 20009 2283 20012
rect 2225 20003 2283 20009
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 7653 20043 7711 20049
rect 7653 20009 7665 20043
rect 7699 20009 7711 20043
rect 7834 20040 7840 20052
rect 7795 20012 7840 20040
rect 7653 20003 7711 20009
rect 1578 19972 1584 19984
rect 1539 19944 1584 19972
rect 1578 19932 1584 19944
rect 1636 19932 1642 19984
rect 7668 19972 7696 20003
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20009 12587 20043
rect 12710 20040 12716 20052
rect 12671 20012 12716 20040
rect 12529 20003 12587 20009
rect 9398 19972 9404 19984
rect 7668 19944 9404 19972
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 12544 19972 12572 20003
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 14645 20043 14703 20049
rect 14645 20009 14657 20043
rect 14691 20009 14703 20043
rect 15010 20040 15016 20052
rect 14971 20012 15016 20040
rect 14645 20003 14703 20009
rect 12802 19972 12808 19984
rect 12544 19944 12808 19972
rect 12802 19932 12808 19944
rect 12860 19972 12866 19984
rect 14660 19972 14688 20003
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 12860 19944 14688 19972
rect 12860 19932 12866 19944
rect 2130 19864 2136 19916
rect 2188 19904 2194 19916
rect 2406 19904 2412 19916
rect 2188 19876 2412 19904
rect 2188 19864 2194 19876
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2590 19864 2596 19916
rect 2648 19904 2654 19916
rect 2777 19907 2835 19913
rect 2777 19904 2789 19907
rect 2648 19876 2789 19904
rect 2648 19864 2654 19876
rect 2777 19873 2789 19876
rect 2823 19873 2835 19907
rect 7558 19904 7564 19916
rect 7519 19876 7564 19904
rect 2777 19867 2835 19873
rect 7558 19864 7564 19876
rect 7616 19864 7622 19916
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 7469 19839 7527 19845
rect 1443 19808 4752 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 2593 19771 2651 19777
rect 2593 19737 2605 19771
rect 2639 19768 2651 19771
rect 3326 19768 3332 19780
rect 2639 19740 3332 19768
rect 2639 19737 2651 19740
rect 2593 19731 2651 19737
rect 3326 19728 3332 19740
rect 3384 19728 3390 19780
rect 4724 19768 4752 19808
rect 7469 19805 7481 19839
rect 7515 19836 7527 19839
rect 8294 19836 8300 19848
rect 7515 19808 8300 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 12342 19836 12348 19848
rect 12303 19808 12348 19836
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 13078 19836 13084 19848
rect 12575 19808 13084 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 14642 19836 14648 19848
rect 14603 19808 14648 19836
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 15746 19836 15752 19848
rect 14875 19808 15752 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 18046 19768 18052 19780
rect 4724 19740 18052 19768
rect 18046 19728 18052 19740
rect 18104 19728 18110 19780
rect 2682 19660 2688 19712
rect 2740 19700 2746 19712
rect 2740 19672 2785 19700
rect 2740 19660 2746 19672
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1397 19499 1455 19505
rect 1397 19465 1409 19499
rect 1443 19496 1455 19499
rect 2682 19496 2688 19508
rect 1443 19468 2688 19496
rect 1443 19465 1455 19468
rect 1397 19459 1455 19465
rect 2682 19456 2688 19468
rect 2740 19456 2746 19508
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 3476 19468 5365 19496
rect 3476 19456 3482 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 5353 19459 5411 19465
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 7745 19499 7803 19505
rect 7745 19496 7757 19499
rect 6963 19468 7757 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7745 19465 7757 19468
rect 7791 19465 7803 19499
rect 7745 19459 7803 19465
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 14875 19468 15669 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 5368 19428 5396 19459
rect 5368 19400 5948 19428
rect 1394 19320 1400 19372
rect 1452 19360 1458 19372
rect 1581 19363 1639 19369
rect 1581 19360 1593 19363
rect 1452 19332 1593 19360
rect 1452 19320 1458 19332
rect 1581 19329 1593 19332
rect 1627 19329 1639 19363
rect 2222 19360 2228 19372
rect 2183 19332 2228 19360
rect 1581 19323 1639 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 2832 19332 3985 19360
rect 2832 19320 2838 19332
rect 3973 19329 3985 19332
rect 4019 19360 4031 19363
rect 4062 19360 4068 19372
rect 4019 19332 4068 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 4240 19363 4298 19369
rect 4240 19329 4252 19363
rect 4286 19360 4298 19363
rect 4286 19332 5856 19360
rect 4286 19329 4298 19332
rect 4240 19323 4298 19329
rect 5828 19224 5856 19332
rect 5920 19292 5948 19400
rect 7098 19388 7104 19440
rect 7156 19428 7162 19440
rect 7156 19400 7880 19428
rect 7156 19388 7162 19400
rect 6549 19363 6607 19369
rect 6549 19329 6561 19363
rect 6595 19360 6607 19363
rect 7561 19363 7619 19369
rect 6595 19332 7512 19360
rect 6595 19329 6607 19332
rect 6549 19323 6607 19329
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 5920 19264 6653 19292
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 7484 19292 7512 19332
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 7650 19360 7656 19372
rect 7607 19332 7656 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 7852 19369 7880 19400
rect 12526 19388 12532 19440
rect 12584 19428 12590 19440
rect 12584 19400 14780 19428
rect 12584 19388 12590 19400
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 8294 19360 8300 19372
rect 7837 19323 7895 19329
rect 7944 19332 8300 19360
rect 7944 19292 7972 19332
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 9398 19360 9404 19372
rect 8588 19332 9404 19360
rect 8386 19292 8392 19304
rect 7484 19264 7972 19292
rect 8347 19264 8392 19292
rect 6641 19255 6699 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 7377 19227 7435 19233
rect 7377 19224 7389 19227
rect 5828 19196 7389 19224
rect 7377 19193 7389 19196
rect 7423 19193 7435 19227
rect 8588 19224 8616 19332
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 12342 19360 12348 19372
rect 11839 19332 12348 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 12342 19320 12348 19332
rect 12400 19360 12406 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12400 19332 12817 19360
rect 12400 19320 12406 19332
rect 12805 19329 12817 19332
rect 12851 19360 12863 19363
rect 14274 19360 14280 19372
rect 12851 19332 14280 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 14274 19320 14280 19332
rect 14332 19360 14338 19372
rect 14461 19363 14519 19369
rect 14461 19360 14473 19363
rect 14332 19332 14473 19360
rect 14332 19320 14338 19332
rect 14461 19329 14473 19332
rect 14507 19360 14519 19363
rect 14642 19360 14648 19372
rect 14507 19332 14648 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 14752 19360 14780 19400
rect 15194 19388 15200 19440
rect 15252 19428 15258 19440
rect 15252 19400 15792 19428
rect 15252 19388 15258 19400
rect 15764 19369 15792 19400
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 14752 19332 15485 19360
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19329 15807 19363
rect 15749 19323 15807 19329
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 7377 19187 7435 19193
rect 8496 19196 8616 19224
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2682 19156 2688 19168
rect 2087 19128 2688 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 8496 19165 8524 19196
rect 6733 19159 6791 19165
rect 6733 19125 6745 19159
rect 6779 19156 6791 19159
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 6779 19128 8493 19156
rect 6779 19125 6791 19128
rect 6733 19119 6791 19125
rect 8481 19125 8493 19128
rect 8527 19125 8539 19159
rect 8662 19156 8668 19168
rect 8623 19128 8668 19156
rect 8481 19119 8539 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 9140 19156 9168 19255
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 9732 19264 11529 19292
rect 9732 19252 9738 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 12894 19292 12900 19304
rect 12855 19264 12900 19292
rect 11517 19255 11575 19261
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 14553 19295 14611 19301
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 16850 19292 16856 19304
rect 14599 19264 16856 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 12250 19184 12256 19236
rect 12308 19224 12314 19236
rect 14568 19224 14596 19255
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 12308 19196 14596 19224
rect 12308 19184 12314 19196
rect 9766 19156 9772 19168
rect 9140 19128 9772 19156
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 12802 19156 12808 19168
rect 12763 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13170 19156 13176 19168
rect 13131 19128 13176 19156
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13722 19116 13728 19168
rect 13780 19156 13786 19168
rect 14461 19159 14519 19165
rect 14461 19156 14473 19159
rect 13780 19128 14473 19156
rect 13780 19116 13786 19128
rect 14461 19125 14473 19128
rect 14507 19125 14519 19159
rect 14461 19119 14519 19125
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15562 19156 15568 19168
rect 15335 19128 15568 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 1912 18924 12434 18952
rect 1912 18912 1918 18924
rect 5445 18887 5503 18893
rect 5445 18853 5457 18887
rect 5491 18884 5503 18887
rect 8386 18884 8392 18896
rect 5491 18856 8392 18884
rect 5491 18853 5503 18856
rect 5445 18847 5503 18853
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 1820 18788 4200 18816
rect 1820 18776 1826 18788
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1412 18680 1440 18711
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2409 18751 2467 18757
rect 2409 18748 2421 18751
rect 2280 18720 2421 18748
rect 2280 18708 2286 18720
rect 2409 18717 2421 18720
rect 2455 18717 2467 18751
rect 4062 18748 4068 18760
rect 4023 18720 4068 18748
rect 2409 18711 2467 18717
rect 4062 18708 4068 18720
rect 4120 18708 4126 18760
rect 4172 18748 4200 18788
rect 5460 18748 5488 18847
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 7742 18776 7748 18828
rect 7800 18816 7806 18828
rect 12406 18816 12434 18924
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13722 18952 13728 18964
rect 12860 18924 13728 18952
rect 12860 18912 12866 18924
rect 13722 18912 13728 18924
rect 13780 18952 13786 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13780 18924 14289 18952
rect 13780 18912 13786 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 16850 18952 16856 18964
rect 16811 18924 16856 18952
rect 14277 18915 14335 18921
rect 16850 18912 16856 18924
rect 16908 18912 16914 18964
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 7800 18788 11100 18816
rect 12406 18788 14381 18816
rect 7800 18776 7806 18788
rect 4172 18720 5488 18748
rect 7561 18751 7619 18757
rect 7561 18717 7573 18751
rect 7607 18748 7619 18751
rect 7650 18748 7656 18760
rect 7607 18720 7656 18748
rect 7607 18717 7619 18720
rect 7561 18711 7619 18717
rect 7650 18708 7656 18720
rect 7708 18708 7714 18760
rect 7837 18751 7895 18757
rect 7837 18717 7849 18751
rect 7883 18748 7895 18751
rect 7926 18748 7932 18760
rect 7883 18720 7932 18748
rect 7883 18717 7895 18720
rect 7837 18711 7895 18717
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9674 18748 9680 18760
rect 9263 18720 9680 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 10962 18748 10968 18760
rect 10192 18720 10968 18748
rect 10192 18708 10198 18720
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 4154 18680 4160 18692
rect 1412 18652 4160 18680
rect 4154 18640 4160 18652
rect 4212 18640 4218 18692
rect 4332 18683 4390 18689
rect 4332 18649 4344 18683
rect 4378 18680 4390 18683
rect 7377 18683 7435 18689
rect 7377 18680 7389 18683
rect 4378 18652 7389 18680
rect 4378 18649 4390 18652
rect 4332 18643 4390 18649
rect 7377 18649 7389 18652
rect 7423 18649 7435 18683
rect 7377 18643 7435 18649
rect 7745 18683 7803 18689
rect 7745 18649 7757 18683
rect 7791 18680 7803 18683
rect 8662 18680 8668 18692
rect 7791 18652 8668 18680
rect 7791 18649 7803 18652
rect 7745 18643 7803 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 1578 18612 1584 18624
rect 1539 18584 1584 18612
rect 1578 18572 1584 18584
rect 1636 18572 1642 18624
rect 2130 18572 2136 18624
rect 2188 18612 2194 18624
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 2188 18584 2237 18612
rect 2188 18572 2194 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 2225 18575 2283 18581
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 9033 18615 9091 18621
rect 9033 18612 9045 18615
rect 8352 18584 9045 18612
rect 8352 18572 8358 18584
rect 9033 18581 9045 18584
rect 9079 18581 9091 18615
rect 11072 18612 11100 18788
rect 14369 18785 14381 18788
rect 14415 18816 14427 18819
rect 14918 18816 14924 18828
rect 14415 18788 14924 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 12989 18751 13047 18757
rect 12989 18748 13001 18751
rect 12584 18720 13001 18748
rect 12584 18708 12590 18720
rect 12989 18717 13001 18720
rect 13035 18717 13047 18751
rect 13170 18748 13176 18760
rect 13131 18720 13176 18748
rect 12989 18711 13047 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 14274 18748 14280 18760
rect 13320 18720 13365 18748
rect 14235 18720 14280 18748
rect 13320 18708 13326 18720
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 11232 18683 11290 18689
rect 11232 18649 11244 18683
rect 11278 18680 11290 18683
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 11278 18652 12817 18680
rect 11278 18649 11290 18652
rect 11232 18643 11290 18649
rect 12805 18649 12817 18652
rect 12851 18649 12863 18683
rect 12805 18643 12863 18649
rect 13446 18640 13452 18692
rect 13504 18680 13510 18692
rect 15488 18680 15516 18711
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 15729 18751 15787 18757
rect 15729 18748 15741 18751
rect 15620 18720 15741 18748
rect 15620 18708 15626 18720
rect 15729 18717 15741 18720
rect 15775 18717 15787 18751
rect 15729 18711 15787 18717
rect 13504 18652 15516 18680
rect 13504 18640 13510 18652
rect 12345 18615 12403 18621
rect 12345 18612 12357 18615
rect 11072 18584 12357 18612
rect 9033 18575 9091 18581
rect 12345 18581 12357 18584
rect 12391 18612 12403 18615
rect 12894 18612 12900 18624
rect 12391 18584 12900 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14645 18615 14703 18621
rect 14645 18581 14657 18615
rect 14691 18612 14703 18615
rect 14734 18612 14740 18624
rect 14691 18584 14740 18612
rect 14691 18581 14703 18584
rect 14645 18575 14703 18581
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 10505 18411 10563 18417
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 10594 18408 10600 18420
rect 10551 18380 10600 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 14918 18408 14924 18420
rect 14879 18380 14924 18408
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 3510 18340 3516 18352
rect 3471 18312 3516 18340
rect 3510 18300 3516 18312
rect 3568 18300 3574 18352
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 15286 18340 15292 18352
rect 4212 18312 15292 18340
rect 4212 18300 4218 18312
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3234 18272 3240 18284
rect 2639 18244 3240 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7708 18244 8033 18272
rect 7708 18232 7714 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 8021 18235 8079 18241
rect 8864 18244 10425 18272
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2740 18176 2789 18204
rect 2740 18164 2746 18176
rect 2777 18173 2789 18176
rect 2823 18173 2835 18207
rect 2777 18167 2835 18173
rect 7558 18164 7564 18216
rect 7616 18204 7622 18216
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 7616 18176 7757 18204
rect 7616 18164 7622 18176
rect 7745 18173 7757 18176
rect 7791 18204 7803 18207
rect 8864 18204 8892 18244
rect 10413 18241 10425 18244
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 12802 18272 12808 18284
rect 11839 18244 12808 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 13808 18275 13866 18281
rect 13808 18241 13820 18275
rect 13854 18272 13866 18275
rect 14366 18272 14372 18284
rect 13854 18244 14372 18272
rect 13854 18241 13866 18244
rect 13808 18235 13866 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 7791 18176 8892 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 9824 18176 11529 18204
rect 9824 18164 9830 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 11517 18167 11575 18173
rect 13464 18176 13553 18204
rect 13464 18080 13492 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 1397 18071 1455 18077
rect 1397 18037 1409 18071
rect 1443 18068 1455 18071
rect 2590 18068 2596 18080
rect 1443 18040 2596 18068
rect 1443 18037 1455 18040
rect 1397 18031 1455 18037
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18068 3847 18071
rect 4982 18068 4988 18080
rect 3835 18040 4988 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 13446 18068 13452 18080
rect 10192 18040 13452 18068
rect 10192 18028 10198 18040
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 18046 17864 18052 17876
rect 18007 17836 18052 17864
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 4062 17688 4068 17740
rect 4120 17728 4126 17740
rect 5905 17731 5963 17737
rect 5905 17728 5917 17731
rect 4120 17700 5917 17728
rect 4120 17688 4126 17700
rect 5905 17697 5917 17700
rect 5951 17697 5963 17731
rect 5905 17691 5963 17697
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 7800 17700 8248 17728
rect 7800 17688 7806 17700
rect 1854 17660 1860 17672
rect 1815 17632 1860 17660
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 2130 17669 2136 17672
rect 2124 17660 2136 17669
rect 2091 17632 2136 17660
rect 2124 17623 2136 17632
rect 2130 17620 2136 17623
rect 2188 17620 2194 17672
rect 2406 17620 2412 17672
rect 2464 17660 2470 17672
rect 2464 17632 2774 17660
rect 2464 17620 2470 17632
rect 2746 17592 2774 17632
rect 7650 17620 7656 17672
rect 7708 17660 7714 17672
rect 8220 17669 8248 17700
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7708 17632 7941 17660
rect 7708 17620 7714 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17629 14611 17663
rect 14826 17660 14832 17672
rect 14787 17632 14832 17660
rect 14553 17623 14611 17629
rect 6172 17595 6230 17601
rect 2746 17564 5856 17592
rect 3234 17524 3240 17536
rect 3195 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 5828 17524 5856 17564
rect 6172 17561 6184 17595
rect 6218 17592 6230 17595
rect 7745 17595 7803 17601
rect 7745 17592 7757 17595
rect 6218 17564 7757 17592
rect 6218 17561 6230 17564
rect 6172 17555 6230 17561
rect 7745 17561 7757 17564
rect 7791 17561 7803 17595
rect 7745 17555 7803 17561
rect 7285 17527 7343 17533
rect 7285 17524 7297 17527
rect 5828 17496 7297 17524
rect 7285 17493 7297 17496
rect 7331 17524 7343 17527
rect 7374 17524 7380 17536
rect 7331 17496 7380 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7708 17496 8125 17524
rect 7708 17484 7714 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 14568 17524 14596 17623
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 16666 17660 16672 17672
rect 16627 17632 16672 17660
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 14734 17592 14740 17604
rect 14695 17564 14740 17592
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 16936 17595 16994 17601
rect 16936 17561 16948 17595
rect 16982 17592 16994 17595
rect 17218 17592 17224 17604
rect 16982 17564 17224 17592
rect 16982 17561 16994 17564
rect 16936 17555 16994 17561
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 15470 17524 15476 17536
rect 14568 17496 15476 17524
rect 8113 17487 8171 17493
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1394 17280 1400 17332
rect 1452 17280 1458 17332
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 7650 17320 7656 17332
rect 7611 17292 7656 17320
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16298 17320 16304 17332
rect 15344 17292 16304 17320
rect 15344 17280 15350 17292
rect 16298 17280 16304 17292
rect 16356 17320 16362 17332
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 16356 17292 18245 17320
rect 16356 17280 16362 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18233 17283 18291 17289
rect 1412 17252 1440 17280
rect 1412 17224 1624 17252
rect 1397 17187 1455 17193
rect 1397 17153 1409 17187
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 1412 17048 1440 17147
rect 1596 17116 1624 17224
rect 7282 17184 7288 17196
rect 7243 17156 7288 17184
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 9766 17184 9772 17196
rect 7432 17156 7477 17184
rect 9727 17156 9772 17184
rect 7432 17144 7438 17156
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10226 17184 10232 17196
rect 10187 17156 10232 17184
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16724 17156 16865 17184
rect 16724 17144 16730 17156
rect 16853 17153 16865 17156
rect 16899 17184 16911 17187
rect 16942 17184 16948 17196
rect 16899 17156 16948 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17120 17187 17178 17193
rect 17120 17153 17132 17187
rect 17166 17184 17178 17187
rect 18138 17184 18144 17196
rect 17166 17156 18144 17184
rect 17166 17153 17178 17156
rect 17120 17147 17178 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 1596 17088 10333 17116
rect 10321 17085 10333 17088
rect 10367 17116 10379 17119
rect 11514 17116 11520 17128
rect 10367 17088 11520 17116
rect 10367 17085 10379 17088
rect 10321 17079 10379 17085
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 13630 17048 13636 17060
rect 1412 17020 13636 17048
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7469 16983 7527 16989
rect 7469 16980 7481 16983
rect 7432 16952 7481 16980
rect 7432 16940 7438 16952
rect 7469 16949 7481 16952
rect 7515 16980 7527 16983
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 7515 16952 9597 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 9585 16949 9597 16952
rect 9631 16980 9643 16983
rect 10318 16980 10324 16992
rect 9631 16952 10324 16980
rect 9631 16949 9643 16952
rect 9585 16943 9643 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16980 10655 16983
rect 12342 16980 12348 16992
rect 10643 16952 12348 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 7374 16776 7380 16788
rect 7335 16748 7380 16776
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 11514 16776 11520 16788
rect 11475 16748 11520 16776
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 16482 16776 16488 16788
rect 16443 16748 16488 16776
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 18138 16776 18144 16788
rect 18099 16748 18144 16776
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 7116 16680 7512 16708
rect 1854 16600 1860 16652
rect 1912 16640 1918 16652
rect 2774 16640 2780 16652
rect 1912 16612 2780 16640
rect 1912 16600 1918 16612
rect 2774 16600 2780 16612
rect 2832 16640 2838 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 2832 16612 4077 16640
rect 2832 16600 2838 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 1412 16504 1440 16535
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 2188 16544 2421 16572
rect 2188 16532 2194 16544
rect 2409 16541 2421 16544
rect 2455 16541 2467 16575
rect 7116 16572 7144 16680
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16609 7435 16643
rect 7377 16603 7435 16609
rect 7282 16572 7288 16584
rect 2409 16535 2467 16541
rect 2746 16544 7144 16572
rect 7243 16544 7288 16572
rect 2746 16504 2774 16544
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 1412 16476 2774 16504
rect 4332 16507 4390 16513
rect 4332 16473 4344 16507
rect 4378 16504 4390 16507
rect 5350 16504 5356 16516
rect 4378 16476 5356 16504
rect 4378 16473 4390 16476
rect 4332 16467 4390 16473
rect 5350 16464 5356 16476
rect 5408 16464 5414 16516
rect 7392 16504 7420 16603
rect 7484 16572 7512 16680
rect 15470 16668 15476 16720
rect 15528 16708 15534 16720
rect 15528 16680 16620 16708
rect 15528 16668 15534 16680
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 16356 16612 16497 16640
rect 16356 16600 16362 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 9306 16572 9312 16584
rect 7484 16544 9312 16572
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10962 16532 10968 16584
rect 11020 16572 11026 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11020 16544 12265 16572
rect 11020 16532 11026 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 12437 16575 12495 16581
rect 12437 16572 12449 16575
rect 12400 16544 12449 16572
rect 12400 16532 12406 16544
rect 12437 16541 12449 16544
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 16206 16572 16212 16584
rect 12575 16544 16212 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16541 16451 16575
rect 16592 16572 16620 16680
rect 17604 16612 17908 16640
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 16592 16544 17417 16572
rect 16393 16535 16451 16541
rect 17405 16541 17417 16544
rect 17451 16572 17463 16575
rect 17604 16572 17632 16612
rect 17451 16544 17632 16572
rect 17681 16575 17739 16581
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17770 16572 17776 16584
rect 17727 16544 17776 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 10226 16504 10232 16516
rect 5460 16476 7420 16504
rect 7576 16476 10232 16504
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2225 16439 2283 16445
rect 2225 16405 2237 16439
rect 2271 16436 2283 16439
rect 2314 16436 2320 16448
rect 2271 16408 2320 16436
rect 2271 16405 2283 16408
rect 2225 16399 2283 16405
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 5460 16445 5488 16476
rect 5445 16439 5503 16445
rect 5445 16436 5457 16439
rect 2556 16408 5457 16436
rect 2556 16396 2562 16408
rect 5445 16405 5457 16408
rect 5491 16405 5503 16439
rect 5445 16399 5503 16405
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7576 16436 7604 16476
rect 7340 16408 7604 16436
rect 7653 16439 7711 16445
rect 7340 16396 7346 16408
rect 7653 16405 7665 16439
rect 7699 16436 7711 16439
rect 7834 16436 7840 16448
rect 7699 16408 7840 16436
rect 7699 16405 7711 16408
rect 7653 16399 7711 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9508 16445 9536 16476
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10404 16507 10462 16513
rect 10404 16473 10416 16507
rect 10450 16504 10462 16507
rect 12069 16507 12127 16513
rect 12069 16504 12081 16507
rect 10450 16476 12081 16504
rect 10450 16473 10462 16476
rect 10404 16467 10462 16473
rect 12069 16473 12081 16476
rect 12115 16473 12127 16507
rect 16408 16504 16436 16535
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 17880 16572 17908 16612
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 17880 16544 18337 16572
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18598 16572 18604 16584
rect 18559 16544 18604 16572
rect 18325 16535 18383 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 16666 16504 16672 16516
rect 16408 16476 16672 16504
rect 12069 16467 12127 16473
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 18509 16507 18567 16513
rect 18509 16504 18521 16507
rect 16776 16476 18521 16504
rect 16776 16445 16804 16476
rect 18509 16473 18521 16476
rect 18555 16473 18567 16507
rect 18509 16467 18567 16473
rect 9493 16439 9551 16445
rect 9493 16405 9505 16439
rect 9539 16405 9551 16439
rect 9493 16399 9551 16405
rect 16761 16439 16819 16445
rect 16761 16405 16773 16439
rect 16807 16405 16819 16439
rect 16761 16399 16819 16405
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 17589 16439 17647 16445
rect 17589 16436 17601 16439
rect 17460 16408 17601 16436
rect 17460 16396 17466 16408
rect 17589 16405 17601 16408
rect 17635 16405 17647 16439
rect 17589 16399 17647 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 1728 16204 2774 16232
rect 1728 16192 1734 16204
rect 2314 16173 2320 16176
rect 2308 16127 2320 16173
rect 2372 16164 2378 16176
rect 2746 16164 2774 16204
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 5408 16204 7481 16232
rect 5408 16192 5414 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 7834 16232 7840 16244
rect 7795 16204 7840 16232
rect 7469 16195 7527 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 17402 16232 17408 16244
rect 17363 16204 17408 16232
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 13446 16164 13452 16176
rect 2372 16136 2408 16164
rect 2746 16136 10456 16164
rect 2314 16124 2320 16127
rect 2372 16124 2378 16136
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1452 16068 1593 16096
rect 1452 16056 1458 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1912 16068 2053 16096
rect 1912 16056 1918 16068
rect 2041 16065 2053 16068
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 6656 16028 6684 16059
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7650 16096 7656 16108
rect 6788 16068 6833 16096
rect 7611 16068 7656 16096
rect 6788 16056 6794 16068
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8018 16096 8024 16108
rect 7975 16068 8024 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8018 16056 8024 16068
rect 8076 16056 8082 16108
rect 10226 16056 10232 16108
rect 10284 16096 10290 16108
rect 10428 16105 10456 16136
rect 11532 16136 13452 16164
rect 11532 16105 11560 16136
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10284 16068 10333 16096
rect 10284 16056 10290 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 7282 16028 7288 16040
rect 6656 16000 7288 16028
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 5810 15960 5816 15972
rect 3344 15932 5816 15960
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 3344 15892 3372 15932
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 7374 15960 7380 15972
rect 6840 15932 7380 15960
rect 1443 15864 3372 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 5074 15892 5080 15904
rect 3476 15864 5080 15892
rect 3476 15852 3482 15864
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 6840 15901 6868 15932
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 10428 15960 10456 16059
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11773 16099 11831 16105
rect 11773 16096 11785 16099
rect 11664 16068 11785 16096
rect 11664 16056 11670 16068
rect 11773 16065 11785 16068
rect 11819 16065 11831 16099
rect 11773 16059 11831 16065
rect 13716 16099 13774 16105
rect 13716 16065 13728 16099
rect 13762 16096 13774 16099
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 13762 16068 15301 16096
rect 13762 16065 13774 16068
rect 13716 16059 13774 16065
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15470 16096 15476 16108
rect 15431 16068 15476 16096
rect 15289 16059 15347 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15654 16096 15660 16108
rect 15615 16068 15660 16096
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 15804 16068 15849 16096
rect 15804 16056 15810 16068
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16724 16068 17049 16096
rect 16724 16056 16730 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 18046 16096 18052 16108
rect 17267 16068 18052 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 13446 16028 13452 16040
rect 13407 16000 13452 16028
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 10428 15932 11284 15960
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15861 6883 15895
rect 7006 15892 7012 15904
rect 6967 15864 7012 15892
rect 6825 15855 6883 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 11146 15892 11152 15904
rect 10735 15864 11152 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11256 15892 11284 15932
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 11256 15864 12909 15892
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 14829 15895 14887 15901
rect 14829 15892 14841 15895
rect 14700 15864 14841 15892
rect 14700 15852 14706 15864
rect 14829 15861 14841 15864
rect 14875 15861 14887 15895
rect 14829 15855 14887 15861
rect 16482 15852 16488 15904
rect 16540 15892 16546 15904
rect 17037 15895 17095 15901
rect 17037 15892 17049 15895
rect 16540 15864 17049 15892
rect 16540 15852 16546 15864
rect 17037 15861 17049 15864
rect 17083 15861 17095 15895
rect 17037 15855 17095 15861
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2240 15660 12434 15688
rect 1486 15580 1492 15632
rect 1544 15620 1550 15632
rect 2240 15620 2268 15660
rect 1544 15592 2268 15620
rect 6641 15623 6699 15629
rect 1544 15580 1550 15592
rect 6641 15589 6653 15623
rect 6687 15620 6699 15623
rect 6730 15620 6736 15632
rect 6687 15592 6736 15620
rect 6687 15589 6699 15592
rect 6641 15583 6699 15589
rect 6730 15580 6736 15592
rect 6788 15580 6794 15632
rect 10781 15623 10839 15629
rect 10781 15589 10793 15623
rect 10827 15620 10839 15623
rect 11606 15620 11612 15632
rect 10827 15592 11612 15620
rect 10827 15589 10839 15592
rect 10781 15583 10839 15589
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 12406 15620 12434 15660
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 14240 15660 14473 15688
rect 14240 15648 14246 15660
rect 14461 15657 14473 15660
rect 14507 15688 14519 15691
rect 14829 15691 14887 15697
rect 14507 15660 14780 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 14642 15620 14648 15632
rect 12406 15592 14648 15620
rect 14642 15580 14648 15592
rect 14700 15580 14706 15632
rect 14752 15620 14780 15660
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 15654 15688 15660 15700
rect 14875 15660 15660 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 17221 15691 17279 15697
rect 17221 15688 17233 15691
rect 16546 15660 17233 15688
rect 16546 15632 16574 15660
rect 17221 15657 17233 15660
rect 17267 15657 17279 15691
rect 17221 15651 17279 15657
rect 16482 15620 16488 15632
rect 14752 15592 16488 15620
rect 16482 15580 16488 15592
rect 16540 15592 16574 15632
rect 16540 15580 16546 15592
rect 2590 15552 2596 15564
rect 2551 15524 2596 15552
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2740 15524 2785 15552
rect 2740 15512 2746 15524
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 7064 15524 7880 15552
rect 7064 15512 7070 15524
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 3418 15484 3424 15496
rect 2547 15456 3424 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 5261 15487 5319 15493
rect 5261 15453 5273 15487
rect 5307 15453 5319 15487
rect 7650 15484 7656 15496
rect 7563 15456 7656 15484
rect 5261 15447 5319 15453
rect 1854 15376 1860 15428
rect 1912 15416 1918 15428
rect 5276 15416 5304 15447
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 7852 15493 7880 15524
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15484 7987 15487
rect 8202 15484 8208 15496
rect 7975 15456 8208 15484
rect 7975 15453 7987 15456
rect 7929 15447 7987 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 10962 15484 10968 15496
rect 10923 15456 10968 15484
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 12158 15484 12164 15496
rect 11287 15456 12164 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 14458 15484 14464 15496
rect 14419 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 14660 15493 14688 15580
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16724 15456 17233 15484
rect 16724 15444 16730 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 17405 15487 17463 15493
rect 17405 15484 17417 15487
rect 17368 15456 17417 15484
rect 17368 15444 17374 15456
rect 17405 15453 17417 15456
rect 17451 15484 17463 15487
rect 17954 15484 17960 15496
rect 17451 15456 17960 15484
rect 17451 15453 17463 15456
rect 17405 15447 17463 15453
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 1912 15388 5304 15416
rect 5528 15419 5586 15425
rect 1912 15376 1918 15388
rect 5528 15385 5540 15419
rect 5574 15416 5586 15419
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 5574 15388 7481 15416
rect 5574 15385 5586 15388
rect 5528 15379 5586 15385
rect 7469 15385 7481 15388
rect 7515 15385 7527 15419
rect 7668 15416 7696 15444
rect 8294 15416 8300 15428
rect 7668 15388 8300 15416
rect 7469 15379 7527 15385
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 1394 15348 1400 15360
rect 1355 15320 1400 15348
rect 1394 15308 1400 15320
rect 1452 15308 1458 15360
rect 17589 15351 17647 15357
rect 17589 15317 17601 15351
rect 17635 15348 17647 15351
rect 17862 15348 17868 15360
rect 17635 15320 17868 15348
rect 17635 15317 17647 15320
rect 17589 15311 17647 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 18012 15116 18613 15144
rect 18012 15104 18018 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 18601 15107 18659 15113
rect 8294 15076 8300 15088
rect 8207 15048 8300 15076
rect 8294 15036 8300 15048
rect 8352 15076 8358 15088
rect 10962 15076 10968 15088
rect 8352 15048 10968 15076
rect 8352 15036 8358 15048
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 15008 1455 15011
rect 1854 15008 1860 15020
rect 1443 14980 1860 15008
rect 1443 14977 1455 14980
rect 1397 14971 1455 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2372 14980 2421 15008
rect 2372 14968 2378 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 7558 15008 7564 15020
rect 7432 14980 7564 15008
rect 7432 14968 7438 14980
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 10060 15017 10088 15048
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7616 14980 8125 15008
rect 7616 14968 7622 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10229 15011 10287 15017
rect 10229 14977 10241 15011
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 12250 15008 12256 15020
rect 10367 14980 12256 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10244 14940 10272 14971
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 14182 15008 14188 15020
rect 14143 14980 14188 15008
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 17494 15017 17500 15020
rect 17488 14971 17500 15017
rect 17552 15008 17558 15020
rect 17552 14980 17588 15008
rect 17494 14968 17500 14971
rect 17552 14968 17558 14980
rect 11238 14940 11244 14952
rect 10244 14912 11244 14940
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 13906 14940 13912 14952
rect 13867 14912 13912 14940
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 17034 14900 17040 14952
rect 17092 14940 17098 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 17092 14912 17233 14940
rect 17092 14900 17098 14912
rect 17221 14909 17233 14912
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 1578 14872 1584 14884
rect 1539 14844 1584 14872
rect 1578 14832 1584 14844
rect 1636 14832 1642 14884
rect 1946 14832 1952 14884
rect 2004 14872 2010 14884
rect 10318 14872 10324 14884
rect 2004 14844 10324 14872
rect 2004 14832 2010 14844
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 2222 14804 2228 14816
rect 2183 14776 2228 14804
rect 2222 14764 2228 14776
rect 2280 14764 2286 14816
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9272 14776 9873 14804
rect 9272 14764 9278 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9861 14767 9919 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 2314 14600 2320 14612
rect 2275 14572 2320 14600
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 4341 14603 4399 14609
rect 4341 14600 4353 14603
rect 2740 14572 4353 14600
rect 2740 14560 2746 14572
rect 4341 14569 4353 14572
rect 4387 14569 4399 14603
rect 10318 14600 10324 14612
rect 10279 14572 10324 14600
rect 4341 14563 4399 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10873 14603 10931 14609
rect 10873 14600 10885 14603
rect 10560 14572 10885 14600
rect 10560 14560 10566 14572
rect 10873 14569 10885 14572
rect 10919 14569 10931 14603
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 10873 14563 10931 14569
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16540 14572 16681 14600
rect 16540 14560 16546 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 17494 14600 17500 14612
rect 17455 14572 17500 14600
rect 16669 14563 16727 14569
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 2590 14492 2596 14544
rect 2648 14532 2654 14544
rect 2648 14504 3004 14532
rect 2648 14492 2654 14504
rect 2976 14476 3004 14504
rect 1394 14424 1400 14476
rect 1452 14464 1458 14476
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 1452 14436 2789 14464
rect 1452 14424 1458 14436
rect 2777 14433 2789 14436
rect 2823 14433 2835 14467
rect 2958 14464 2964 14476
rect 2919 14436 2964 14464
rect 2777 14427 2835 14433
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 5810 14464 5816 14476
rect 5771 14436 5816 14464
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14464 6055 14467
rect 6270 14464 6276 14476
rect 6043 14436 6276 14464
rect 6043 14433 6055 14436
rect 5997 14427 6055 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 10336 14464 10364 14560
rect 10965 14467 11023 14473
rect 10965 14464 10977 14467
rect 10336 14436 10977 14464
rect 10965 14433 10977 14436
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 15470 14464 15476 14476
rect 13587 14436 15476 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 15470 14424 15476 14436
rect 15528 14464 15534 14476
rect 15528 14436 17724 14464
rect 15528 14424 15534 14436
rect 1578 14396 1584 14408
rect 1539 14368 1584 14396
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9214 14405 9220 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8812 14368 8953 14396
rect 8812 14356 8818 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 9208 14396 9220 14405
rect 9175 14368 9220 14396
rect 8941 14359 8999 14365
rect 9208 14359 9220 14368
rect 9214 14356 9220 14359
rect 9272 14356 9278 14408
rect 10870 14396 10876 14408
rect 10831 14368 10876 14396
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 12952 14368 14105 14396
rect 12952 14356 12958 14368
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14274 14396 14280 14408
rect 14139 14368 14280 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14458 14396 14464 14408
rect 14415 14368 14464 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14458 14356 14464 14368
rect 14516 14396 14522 14408
rect 16666 14396 16672 14408
rect 14516 14368 16672 14396
rect 14516 14356 14522 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16850 14396 16856 14408
rect 16811 14368 16856 14396
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17696 14405 17724 14436
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14365 17739 14399
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 17681 14359 17739 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14396 18015 14399
rect 18230 14396 18236 14408
rect 18003 14368 18236 14396
rect 18003 14365 18015 14368
rect 17957 14359 18015 14365
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 1412 14300 3924 14328
rect 1412 14269 1440 14300
rect 1397 14263 1455 14269
rect 1397 14229 1409 14263
rect 1443 14229 1455 14263
rect 2682 14260 2688 14272
rect 2643 14232 2688 14260
rect 1397 14223 1455 14229
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 3896 14260 3924 14300
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 4028 14300 4261 14328
rect 4028 14288 4034 14300
rect 4249 14297 4261 14300
rect 4295 14297 4307 14331
rect 13354 14328 13360 14340
rect 13315 14300 13360 14328
rect 4249 14291 4307 14297
rect 13354 14288 13360 14300
rect 13412 14288 13418 14340
rect 4614 14260 4620 14272
rect 3896 14232 4620 14260
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 5350 14260 5356 14272
rect 5311 14232 5356 14260
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5718 14260 5724 14272
rect 5679 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 16850 14260 16856 14272
rect 13688 14232 16856 14260
rect 13688 14220 13694 14232
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17037 14263 17095 14269
rect 17037 14229 17049 14263
rect 17083 14260 17095 14263
rect 17218 14260 17224 14272
rect 17083 14232 17224 14260
rect 17083 14229 17095 14232
rect 17037 14223 17095 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2096 14028 2360 14056
rect 2096 14016 2102 14028
rect 2222 13997 2228 14000
rect 2216 13988 2228 13997
rect 2183 13960 2228 13988
rect 2216 13951 2228 13960
rect 2222 13948 2228 13951
rect 2280 13948 2286 14000
rect 2332 13988 2360 14028
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 3329 14059 3387 14065
rect 3329 14056 3341 14059
rect 2740 14028 3341 14056
rect 2740 14016 2746 14028
rect 3329 14025 3341 14028
rect 3375 14056 3387 14059
rect 8478 14056 8484 14068
rect 3375 14028 8484 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13446 14056 13452 14068
rect 12768 14028 13452 14056
rect 12768 14016 12774 14028
rect 13446 14016 13452 14028
rect 13504 14056 13510 14068
rect 13504 14028 16574 14056
rect 13504 14016 13510 14028
rect 2332 13960 14780 13988
rect 1762 13880 1768 13932
rect 1820 13920 1826 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1820 13892 1961 13920
rect 1820 13880 1826 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 3970 13920 3976 13932
rect 3927 13892 3976 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5408 13892 5733 13920
rect 5408 13880 5414 13892
rect 5721 13889 5733 13892
rect 5767 13889 5779 13923
rect 12710 13920 12716 13932
rect 12671 13892 12716 13920
rect 5721 13883 5779 13889
rect 12710 13880 12716 13892
rect 12768 13880 12774 13932
rect 12980 13923 13038 13929
rect 12980 13889 12992 13923
rect 13026 13920 13038 13923
rect 14090 13920 14096 13932
rect 13026 13892 14096 13920
rect 13026 13889 13038 13892
rect 12980 13883 13038 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 2958 13812 2964 13864
rect 3016 13852 3022 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 3016 13824 4077 13852
rect 3016 13812 3022 13824
rect 4065 13821 4077 13824
rect 4111 13852 4123 13855
rect 6270 13852 6276 13864
rect 4111 13824 6276 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 9824 13824 10149 13852
rect 9824 13812 9830 13824
rect 10137 13821 10149 13824
rect 10183 13852 10195 13855
rect 10226 13852 10232 13864
rect 10183 13824 10232 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10502 13852 10508 13864
rect 10459 13824 10508 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13784 14151 13787
rect 14200 13784 14228 13960
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14752 13929 14780 13960
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 14332 13892 14657 13920
rect 14332 13880 14338 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14139 13756 14228 13784
rect 16546 13852 16574 14028
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 16908 14028 18061 14056
rect 16908 14016 16914 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 16942 13929 16948 13932
rect 16936 13883 16948 13929
rect 17000 13920 17006 13932
rect 17000 13892 17036 13920
rect 16942 13880 16948 13883
rect 17000 13880 17006 13892
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16546 13824 16681 13852
rect 14139 13753 14151 13756
rect 14093 13747 14151 13753
rect 5537 13719 5595 13725
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 5810 13716 5816 13728
rect 5583 13688 5816 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14645 13719 14703 13725
rect 14645 13716 14657 13719
rect 13964 13688 14657 13716
rect 13964 13676 13970 13688
rect 14645 13685 14657 13688
rect 14691 13685 14703 13719
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 14645 13679 14703 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 16546 13716 16574 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 16850 13716 16856 13728
rect 16546 13688 16856 13716
rect 16850 13676 16856 13688
rect 16908 13716 16914 13728
rect 17034 13716 17040 13728
rect 16908 13688 17040 13716
rect 16908 13676 16914 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 2406 13472 2412 13524
rect 2464 13512 2470 13524
rect 5626 13512 5632 13524
rect 2464 13484 5632 13512
rect 2464 13472 2470 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 6822 13512 6828 13524
rect 5776 13484 6828 13512
rect 5776 13472 5782 13484
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 10502 13512 10508 13524
rect 9539 13484 10508 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 14090 13512 14096 13524
rect 14051 13484 14096 13512
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 16853 13515 16911 13521
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 16942 13512 16948 13524
rect 16899 13484 16948 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 1412 13348 5580 13376
rect 1412 13317 1440 13348
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3568 13280 3801 13308
rect 3568 13268 3574 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13277 5503 13311
rect 5445 13271 5503 13277
rect 3970 13172 3976 13184
rect 3931 13144 3976 13172
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 5460 13172 5488 13271
rect 5552 13240 5580 13348
rect 9324 13348 10456 13376
rect 5718 13317 5724 13320
rect 5701 13311 5724 13317
rect 5701 13277 5713 13311
rect 5701 13271 5724 13277
rect 5718 13268 5724 13271
rect 5776 13268 5782 13320
rect 9324 13317 9352 13348
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9456 13280 9501 13308
rect 9456 13268 9462 13280
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 10042 13308 10048 13320
rect 9732 13280 10048 13308
rect 9732 13268 9738 13280
rect 10042 13268 10048 13280
rect 10100 13308 10106 13320
rect 10428 13317 10456 13348
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 10560 13348 12725 13376
rect 10560 13336 10566 13348
rect 12713 13345 12725 13348
rect 12759 13376 12771 13379
rect 13906 13376 13912 13388
rect 12759 13348 13912 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 10100 13280 10149 13308
rect 10100 13268 10106 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13308 10471 13311
rect 10870 13308 10876 13320
rect 10459 13280 10876 13308
rect 10459 13277 10471 13280
rect 10413 13271 10471 13277
rect 10870 13268 10876 13280
rect 10928 13308 10934 13320
rect 12894 13308 12900 13320
rect 10928 13280 12900 13308
rect 10928 13268 10934 13280
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13170 13308 13176 13320
rect 13035 13280 13176 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 13722 13308 13728 13320
rect 13412 13280 13728 13308
rect 13412 13268 13418 13280
rect 13722 13268 13728 13280
rect 13780 13308 13786 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 13780 13280 14289 13308
rect 13780 13268 13786 13280
rect 14277 13277 14289 13280
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 15562 13308 15568 13320
rect 14599 13280 15568 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 15562 13268 15568 13280
rect 15620 13268 15626 13320
rect 17037 13311 17095 13317
rect 17037 13277 17049 13311
rect 17083 13277 17095 13311
rect 17218 13308 17224 13320
rect 17179 13280 17224 13308
rect 17037 13271 17095 13277
rect 14461 13243 14519 13249
rect 5552 13212 14412 13240
rect 5534 13172 5540 13184
rect 5460 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 5626 13132 5632 13184
rect 5684 13172 5690 13184
rect 9398 13172 9404 13184
rect 5684 13144 9404 13172
rect 5684 13132 5690 13144
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 10502 13172 10508 13184
rect 9723 13144 10508 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 14384 13172 14412 13212
rect 14461 13209 14473 13243
rect 14507 13240 14519 13243
rect 15010 13240 15016 13252
rect 14507 13212 15016 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 17052 13240 17080 13271
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17494 13308 17500 13320
rect 17359 13280 17500 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17126 13240 17132 13252
rect 17052 13212 17132 13240
rect 17126 13200 17132 13212
rect 17184 13200 17190 13252
rect 15838 13172 15844 13184
rect 14384 13144 15844 13172
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 10137 12971 10195 12977
rect 10137 12968 10149 12971
rect 9456 12940 10149 12968
rect 9456 12928 9462 12940
rect 10137 12937 10149 12940
rect 10183 12937 10195 12971
rect 10137 12931 10195 12937
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 15896 12940 18429 12968
rect 15896 12928 15902 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 12342 12900 12348 12912
rect 1412 12872 12348 12900
rect 1412 12841 1440 12872
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 14642 12900 14648 12912
rect 14555 12872 14648 12900
rect 14642 12860 14648 12872
rect 14700 12900 14706 12912
rect 17126 12900 17132 12912
rect 14700 12872 17132 12900
rect 14700 12860 14706 12872
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 1397 12795 1455 12801
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 5718 12832 5724 12844
rect 4571 12804 5724 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6733 12835 6791 12841
rect 5859 12804 6408 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 6270 12764 6276 12776
rect 4847 12736 6276 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4614 12628 4620 12640
rect 4203 12600 4620 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5626 12628 5632 12640
rect 5587 12600 5632 12628
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6380 12637 6408 12804
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 7650 12832 7656 12844
rect 6779 12804 7656 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9024 12835 9082 12841
rect 9024 12801 9036 12835
rect 9070 12832 9082 12835
rect 10134 12832 10140 12844
rect 9070 12804 10140 12832
rect 9070 12801 9082 12804
rect 9024 12795 9082 12801
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10244 12804 10793 12832
rect 6454 12724 6460 12776
rect 6512 12764 6518 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6512 12736 6837 12764
rect 6512 12724 6518 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 6546 12656 6552 12708
rect 6604 12696 6610 12708
rect 6932 12696 6960 12727
rect 6604 12668 6960 12696
rect 6604 12656 6610 12668
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12597 6423 12631
rect 6365 12591 6423 12597
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 10244 12628 10272 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12952 12804 13093 12832
rect 12952 12792 12958 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13722 12696 13728 12708
rect 12406 12668 13728 12696
rect 7432 12600 10272 12628
rect 7432 12588 7438 12600
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10376 12600 10885 12628
rect 10376 12588 10382 12600
rect 10873 12597 10885 12600
rect 10919 12628 10931 12631
rect 12406 12628 12434 12668
rect 13722 12656 13728 12668
rect 13780 12696 13786 12708
rect 14476 12696 14504 12795
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15344 12804 15761 12832
rect 15344 12792 15350 12804
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 15896 12804 15941 12832
rect 15896 12792 15902 12804
rect 16942 12792 16948 12844
rect 17000 12832 17006 12844
rect 17293 12835 17351 12841
rect 17293 12832 17305 12835
rect 17000 12804 17305 12832
rect 17000 12792 17006 12804
rect 17293 12801 17305 12804
rect 17339 12801 17351 12835
rect 17293 12795 17351 12801
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16908 12736 17049 12764
rect 16908 12724 16914 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 13780 12668 14504 12696
rect 13780 12656 13786 12668
rect 10919 12600 12434 12628
rect 10919 12597 10931 12600
rect 10873 12591 10931 12597
rect 15378 12588 15384 12640
rect 15436 12628 15442 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15436 12600 15761 12628
rect 15436 12588 15442 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 17310 12628 17316 12640
rect 16163 12600 17316 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2406 12424 2412 12436
rect 2271 12396 2412 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 6454 12424 6460 12436
rect 2746 12396 6460 12424
rect 1397 12359 1455 12365
rect 1397 12325 1409 12359
rect 1443 12356 1455 12359
rect 2746 12356 2774 12396
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12400 12396 13093 12424
rect 12400 12384 12406 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 1443 12328 2774 12356
rect 1443 12325 1455 12328
rect 1397 12319 1455 12325
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2648 12260 2789 12288
rect 2648 12248 2654 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 13096 12288 13124 12387
rect 13170 12384 13176 12436
rect 13228 12424 13234 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13228 12396 14289 12424
rect 13228 12384 13234 12396
rect 14277 12393 14289 12396
rect 14323 12424 14335 12427
rect 15378 12424 15384 12436
rect 14323 12396 15384 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 16942 12424 16948 12436
rect 16903 12396 16948 12424
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 13262 12316 13268 12368
rect 13320 12356 13326 12368
rect 13446 12356 13452 12368
rect 13320 12328 13452 12356
rect 13320 12316 13326 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 2777 12251 2835 12257
rect 10612 12260 11836 12288
rect 13096 12260 14197 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1452 12192 1593 12220
rect 1452 12180 1458 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4614 12220 4620 12232
rect 4571 12192 4620 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 6144 12192 6285 12220
rect 6144 12180 6150 12192
rect 6273 12189 6285 12192
rect 6319 12220 6331 12223
rect 8754 12220 8760 12232
rect 6319 12192 8760 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10612 12229 10640 12260
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 11698 12220 11704 12232
rect 11659 12192 11704 12220
rect 10597 12183 10655 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11808 12220 11836 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 11808 12192 12664 12220
rect 2593 12155 2651 12161
rect 2593 12121 2605 12155
rect 2639 12152 2651 12155
rect 3234 12152 3240 12164
rect 2639 12124 3240 12152
rect 2639 12121 2651 12124
rect 2593 12115 2651 12121
rect 3234 12112 3240 12124
rect 3292 12112 3298 12164
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 6518 12155 6576 12161
rect 6518 12152 6530 12155
rect 5684 12124 6530 12152
rect 5684 12112 5690 12124
rect 6518 12121 6530 12124
rect 6564 12121 6576 12155
rect 6518 12115 6576 12121
rect 11968 12155 12026 12161
rect 11968 12121 11980 12155
rect 12014 12152 12026 12155
rect 12636 12152 12664 12192
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13354 12220 13360 12232
rect 12768 12192 13360 12220
rect 12768 12180 12774 12192
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13412 12192 14105 12220
rect 13412 12180 13418 12192
rect 14093 12189 14105 12192
rect 14139 12220 14151 12223
rect 15286 12220 15292 12232
rect 14139 12192 15292 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 17126 12220 17132 12232
rect 17087 12192 17132 12220
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 17310 12220 17316 12232
rect 17271 12192 17316 12220
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 17460 12192 17505 12220
rect 17460 12180 17466 12192
rect 16666 12152 16672 12164
rect 12014 12124 12434 12152
rect 12636 12124 16672 12152
rect 12014 12121 12026 12124
rect 11968 12115 12026 12121
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 4338 12084 4344 12096
rect 2740 12056 2785 12084
rect 4299 12056 4344 12084
rect 2740 12044 2746 12056
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 12406 12084 12434 12124
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 12526 12084 12532 12096
rect 12406 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 13688 12056 14473 12084
rect 13688 12044 13694 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 1912 11852 7604 11880
rect 1912 11840 1918 11852
rect 2124 11815 2182 11821
rect 2124 11781 2136 11815
rect 2170 11812 2182 11815
rect 2222 11812 2228 11824
rect 2170 11784 2228 11812
rect 2170 11781 2182 11784
rect 2124 11775 2182 11781
rect 2222 11772 2228 11784
rect 2280 11772 2286 11824
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4678 11815 4736 11821
rect 4678 11812 4690 11815
rect 4396 11784 4690 11812
rect 4396 11772 4402 11784
rect 4678 11781 4690 11784
rect 4724 11781 4736 11815
rect 4678 11775 4736 11781
rect 1762 11704 1768 11756
rect 1820 11744 1826 11756
rect 1857 11747 1915 11753
rect 1857 11744 1869 11747
rect 1820 11716 1869 11744
rect 1820 11704 1826 11716
rect 1857 11713 1869 11716
rect 1903 11744 1915 11747
rect 2498 11744 2504 11756
rect 1903 11716 2504 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 2498 11704 2504 11716
rect 2556 11744 2562 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 2556 11716 4445 11744
rect 2556 11704 2562 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 5534 11744 5540 11756
rect 4479 11716 5540 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 5534 11704 5540 11716
rect 5592 11744 5598 11756
rect 6086 11744 6092 11756
rect 5592 11716 6092 11744
rect 5592 11704 5598 11716
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 7576 11676 7604 11852
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 12584 11852 13277 11880
rect 12584 11840 12590 11852
rect 13265 11849 13277 11852
rect 13311 11849 13323 11883
rect 13630 11880 13636 11892
rect 13591 11852 13636 11880
rect 13265 11843 13323 11849
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 11977 11815 12035 11821
rect 11977 11812 11989 11815
rect 10376 11784 11989 11812
rect 10376 11772 10382 11784
rect 11977 11781 11989 11784
rect 12023 11781 12035 11815
rect 14642 11812 14648 11824
rect 11977 11775 12035 11781
rect 13464 11784 14648 11812
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 7708 11716 8309 11744
rect 7708 11704 7714 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8662 11744 8668 11756
rect 8527 11716 8668 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 13354 11744 13360 11756
rect 9364 11716 13360 11744
rect 9364 11704 9370 11716
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 13464 11753 13492 11784
rect 14642 11772 14648 11784
rect 14700 11772 14706 11824
rect 16758 11812 16764 11824
rect 15120 11784 16764 11812
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 15120 11744 15148 11784
rect 16758 11772 16764 11784
rect 16816 11772 16822 11824
rect 15286 11744 15292 11756
rect 13771 11716 15148 11744
rect 15247 11716 15292 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 15286 11704 15292 11716
rect 15344 11744 15350 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 15344 11716 16957 11744
rect 15344 11704 15350 11716
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 7576 11648 15393 11676
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 15930 11676 15936 11688
rect 15427 11648 15936 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 17037 11679 17095 11685
rect 17037 11645 17049 11679
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 9766 11608 9772 11620
rect 6880 11580 9772 11608
rect 6880 11568 6886 11580
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 17052 11608 17080 11639
rect 18690 11608 18696 11620
rect 15304 11580 18696 11608
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 5810 11540 5816 11552
rect 5771 11512 5816 11540
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 8665 11543 8723 11549
rect 8665 11509 8677 11543
rect 8711 11540 8723 11543
rect 11238 11540 11244 11552
rect 8711 11512 11244 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11974 11500 11980 11552
rect 12032 11540 12038 11552
rect 12069 11543 12127 11549
rect 12069 11540 12081 11543
rect 12032 11512 12081 11540
rect 12032 11500 12038 11512
rect 12069 11509 12081 11512
rect 12115 11509 12127 11543
rect 12069 11503 12127 11509
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 15304 11540 15332 11580
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 13412 11512 15332 11540
rect 13412 11500 13418 11512
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 15436 11512 15485 11540
rect 15436 11500 15442 11512
rect 15473 11509 15485 11512
rect 15519 11540 15531 11543
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 15519 11512 16957 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17313 11543 17371 11549
rect 17313 11509 17325 11543
rect 17359 11540 17371 11543
rect 17862 11540 17868 11552
rect 17359 11512 17868 11540
rect 17359 11509 17371 11512
rect 17313 11503 17371 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 13170 11336 13176 11348
rect 12851 11308 13176 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 15930 11336 15936 11348
rect 15891 11308 15936 11336
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 1578 11268 1584 11280
rect 1539 11240 1584 11268
rect 1578 11228 1584 11240
rect 1636 11228 1642 11280
rect 2133 11271 2191 11277
rect 2133 11237 2145 11271
rect 2179 11268 2191 11271
rect 3050 11268 3056 11280
rect 2179 11240 3056 11268
rect 2179 11237 2191 11240
rect 2133 11231 2191 11237
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 3234 11228 3240 11280
rect 3292 11268 3298 11280
rect 3292 11240 8984 11268
rect 3292 11228 3298 11240
rect 8956 11209 8984 11240
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12526 11268 12532 11280
rect 11756 11240 12532 11268
rect 11756 11228 11762 11240
rect 12526 11228 12532 11240
rect 12584 11268 12590 11280
rect 12584 11240 14596 11268
rect 12584 11228 12590 11240
rect 8941 11203 8999 11209
rect 1412 11172 5764 11200
rect 1412 11141 1440 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2774 11132 2780 11144
rect 2363 11104 2780 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 5736 11064 5764 11172
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9646 11172 9996 11200
rect 5810 11092 5816 11144
rect 5868 11132 5874 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 5868 11104 8033 11132
rect 5868 11092 5874 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8662 11132 8668 11144
rect 8251 11104 8668 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8662 11092 8668 11104
rect 8720 11132 8726 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8720 11104 9137 11132
rect 8720 11092 8726 11104
rect 9039 11100 9076 11104
rect 9125 11101 9137 11104
rect 9171 11132 9183 11135
rect 9646 11132 9674 11172
rect 9171 11104 9674 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 9968 11141 9996 11172
rect 12406 11172 12848 11200
rect 9953 11135 10011 11141
rect 9824 11104 9869 11132
rect 9824 11092 9830 11104
rect 9953 11101 9965 11135
rect 9999 11101 10011 11135
rect 12406 11132 12434 11172
rect 12820 11144 12848 11172
rect 12618 11132 12624 11144
rect 9953 11095 10011 11101
rect 10060 11104 12434 11132
rect 12579 11104 12624 11132
rect 9306 11064 9312 11076
rect 5736 11036 9168 11064
rect 9267 11036 9312 11064
rect 8386 10996 8392 11008
rect 8347 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 9140 10996 9168 11036
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 10060 10996 10088 11104
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 12802 11132 12808 11144
rect 12763 11104 12808 11132
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 14568 11141 14596 11240
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 16850 11132 16856 11144
rect 14599 11104 16856 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 16850 11092 16856 11104
rect 16908 11132 16914 11144
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 16908 11104 17325 11132
rect 16908 11092 16914 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 10137 11067 10195 11073
rect 10137 11033 10149 11067
rect 10183 11064 10195 11067
rect 10870 11064 10876 11076
rect 10183 11036 10876 11064
rect 10183 11033 10195 11036
rect 10137 11027 10195 11033
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 14820 11067 14878 11073
rect 14820 11033 14832 11067
rect 14866 11064 14878 11067
rect 15286 11064 15292 11076
rect 14866 11036 15292 11064
rect 14866 11033 14878 11036
rect 14820 11027 14878 11033
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 17586 11073 17592 11076
rect 17580 11027 17592 11073
rect 17644 11064 17650 11076
rect 17644 11036 17680 11064
rect 17586 11024 17592 11027
rect 17644 11024 17650 11036
rect 9140 10968 10088 10996
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12989 10999 13047 11005
rect 12989 10996 13001 10999
rect 12492 10968 13001 10996
rect 12492 10956 12498 10968
rect 12989 10965 13001 10968
rect 13035 10965 13047 10999
rect 12989 10959 13047 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 2682 10792 2688 10804
rect 1443 10764 2688 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 12860 10764 12909 10792
rect 12860 10752 12866 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 12897 10755 12955 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15654 10792 15660 10804
rect 15615 10764 15660 10792
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17586 10792 17592 10804
rect 17543 10764 17592 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 17126 10724 17132 10736
rect 15488 10696 17132 10724
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1452 10628 1593 10656
rect 1452 10616 1458 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3878 10656 3884 10668
rect 3007 10628 3884 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 8478 10656 8484 10668
rect 8439 10628 8484 10656
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 11784 10659 11842 10665
rect 11784 10625 11796 10659
rect 11830 10656 11842 10659
rect 12066 10656 12072 10668
rect 11830 10628 12072 10656
rect 11830 10625 11842 10628
rect 11784 10619 11842 10625
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 15488 10665 15516 10696
rect 17126 10684 17132 10696
rect 17184 10724 17190 10736
rect 17184 10696 17724 10724
rect 17184 10684 17190 10696
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 16574 10656 16580 10668
rect 15795 10628 16580 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 17696 10665 17724 10696
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17957 10659 18015 10665
rect 17957 10625 17969 10659
rect 18003 10656 18015 10659
rect 19334 10656 19340 10668
rect 18003 10628 19340 10656
rect 18003 10625 18015 10628
rect 17957 10619 18015 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 3234 10588 3240 10600
rect 3195 10560 3240 10588
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11480 10560 11529 10588
rect 11480 10548 11486 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10452 2651 10455
rect 2866 10452 2872 10464
rect 2639 10424 2872 10452
rect 2639 10421 2651 10424
rect 2593 10415 2651 10421
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 9582 10452 9588 10464
rect 8895 10424 9588 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10217 5319 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5261 10211 5319 10217
rect 5276 10180 5304 10211
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8662 10248 8668 10260
rect 7975 10220 8668 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 12066 10248 12072 10260
rect 12027 10220 12072 10248
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 5626 10180 5632 10192
rect 5276 10152 5632 10180
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 5132 10084 5181 10112
rect 5132 10072 5138 10084
rect 5169 10081 5181 10084
rect 5215 10112 5227 10115
rect 5350 10112 5356 10124
rect 5215 10084 5356 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3326 10004 3332 10056
rect 3384 10044 3390 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 3384 10016 4997 10044
rect 3384 10004 3390 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5718 10044 5724 10056
rect 5307 10016 5724 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6086 10044 6092 10056
rect 5999 10016 6092 10044
rect 6086 10004 6092 10016
rect 6144 10044 6150 10056
rect 8110 10044 8116 10056
rect 6144 10016 6592 10044
rect 8071 10016 8116 10044
rect 6144 10004 6150 10016
rect 6564 9988 6592 10016
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12032 10016 12265 10044
rect 12032 10004 12038 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 13998 10044 14004 10056
rect 12575 10016 14004 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 6362 9985 6368 9988
rect 6356 9939 6368 9985
rect 6420 9976 6426 9988
rect 6420 9948 6456 9976
rect 6362 9936 6368 9939
rect 6420 9936 6426 9948
rect 6546 9936 6552 9988
rect 6604 9936 6610 9988
rect 2685 9911 2743 9917
rect 2685 9877 2697 9911
rect 2731 9908 2743 9911
rect 2774 9908 2780 9920
rect 2731 9880 2780 9908
rect 2731 9877 2743 9880
rect 2685 9871 2743 9877
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 8846 9908 8852 9920
rect 7515 9880 8852 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12492 9880 12537 9908
rect 12492 9868 12498 9880
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 6362 9704 6368 9716
rect 6323 9676 6368 9704
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 8941 9707 8999 9713
rect 8941 9673 8953 9707
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 2774 9645 2780 9648
rect 2768 9599 2780 9645
rect 2832 9636 2838 9648
rect 2832 9608 2868 9636
rect 2774 9596 2780 9599
rect 2832 9596 2838 9608
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 6086 9568 6092 9580
rect 1443 9540 6092 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6236 9540 6561 9568
rect 6236 9528 6242 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 8956 9568 8984 9667
rect 19242 9636 19248 9648
rect 12406 9608 19248 9636
rect 10042 9568 10048 9580
rect 8076 9540 8616 9568
rect 8956 9540 10048 9568
rect 8076 9528 8082 9540
rect 2498 9500 2504 9512
rect 2459 9472 2504 9500
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 7892 9472 8493 9500
rect 7892 9460 7898 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8588 9500 8616 9540
rect 10042 9528 10048 9540
rect 10100 9528 10106 9580
rect 12406 9568 12434 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 15746 9568 15752 9580
rect 10152 9540 12434 9568
rect 15707 9540 15752 9568
rect 10152 9500 10180 9540
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 16925 9571 16983 9577
rect 16925 9568 16937 9571
rect 16080 9540 16937 9568
rect 16080 9528 16086 9540
rect 16925 9537 16937 9540
rect 16971 9537 16983 9571
rect 16925 9531 16983 9537
rect 10318 9500 10324 9512
rect 8588 9472 10180 9500
rect 10279 9472 10324 9500
rect 8481 9463 8539 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 15841 9503 15899 9509
rect 15841 9500 15853 9503
rect 10428 9472 15853 9500
rect 8846 9432 8852 9444
rect 8807 9404 8852 9432
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 3878 9364 3884 9376
rect 3839 9336 3884 9364
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 10428 9364 10456 9472
rect 15841 9469 15853 9472
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9500 15991 9503
rect 16482 9500 16488 9512
rect 15979 9472 16488 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 11422 9392 11428 9444
rect 11480 9432 11486 9444
rect 12526 9432 12532 9444
rect 11480 9404 12532 9432
rect 11480 9392 11486 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 5868 9336 10456 9364
rect 15381 9367 15439 9373
rect 5868 9324 5874 9336
rect 15381 9333 15393 9367
rect 15427 9364 15439 9367
rect 16114 9364 16120 9376
rect 15427 9336 16120 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16684 9364 16712 9463
rect 16850 9364 16856 9376
rect 16684 9336 16856 9364
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 18046 9364 18052 9376
rect 18007 9336 18052 9364
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 5810 9160 5816 9172
rect 1728 9132 5816 9160
rect 1728 9120 1734 9132
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 5994 9160 6000 9172
rect 5955 9132 6000 9160
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 10962 9160 10968 9172
rect 9692 9132 10968 9160
rect 1397 9095 1455 9101
rect 1397 9061 1409 9095
rect 1443 9092 1455 9095
rect 2958 9092 2964 9104
rect 1443 9064 2964 9092
rect 1443 9061 1455 9064
rect 1397 9055 1455 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 3234 9092 3240 9104
rect 3195 9064 3240 9092
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 5626 9092 5632 9104
rect 5587 9064 5632 9092
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 9692 9092 9720 9132
rect 10962 9120 10968 9132
rect 11020 9160 11026 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11020 9132 11989 9160
rect 11020 9120 11026 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16022 9160 16028 9172
rect 15979 9132 16028 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 19242 9160 19248 9172
rect 19203 9132 19248 9160
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 6144 9064 9720 9092
rect 6144 9052 6150 9064
rect 12250 9052 12256 9104
rect 12308 9092 12314 9104
rect 17681 9095 17739 9101
rect 17681 9092 17693 9095
rect 12308 9064 17693 9092
rect 12308 9052 12314 9064
rect 17681 9061 17693 9064
rect 17727 9061 17739 9095
rect 17681 9055 17739 9061
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2774 8956 2780 8968
rect 2271 8928 2780 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2774 8916 2780 8928
rect 2832 8916 2838 8968
rect 3050 8956 3056 8968
rect 2963 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8956 3114 8968
rect 3510 8956 3516 8968
rect 3108 8928 3516 8956
rect 3108 8916 3114 8928
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 5644 8956 5672 9052
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 7742 9024 7748 9036
rect 7607 8996 7748 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 7742 8984 7748 8996
rect 7800 9024 7806 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 7800 8996 9137 9024
rect 7800 8984 7806 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10226 9024 10232 9036
rect 10091 8996 10232 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 7834 8956 7840 8968
rect 5644 8928 7840 8956
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 8720 8928 9229 8956
rect 8720 8916 8726 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8956 10655 8959
rect 11422 8956 11428 8968
rect 10643 8928 11428 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 10612 8888 10640 8919
rect 11422 8916 11428 8928
rect 11480 8916 11486 8968
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 16114 8956 16120 8968
rect 16075 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 17862 8956 17868 8968
rect 17823 8928 17868 8956
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 19150 8956 19156 8968
rect 18187 8928 19156 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19426 8956 19432 8968
rect 19387 8928 19432 8956
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20622 8956 20628 8968
rect 19751 8928 20628 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 10100 8860 10640 8888
rect 10864 8891 10922 8897
rect 10100 8848 10106 8860
rect 10864 8857 10876 8891
rect 10910 8888 10922 8891
rect 11514 8888 11520 8900
rect 10910 8860 11520 8888
rect 10910 8857 10922 8860
rect 10864 8851 10922 8857
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 19058 8888 19064 8900
rect 12216 8860 19064 8888
rect 12216 8848 12222 8860
rect 19058 8848 19064 8860
rect 19116 8848 19122 8900
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 13170 8820 13176 8832
rect 13131 8792 13176 8820
rect 5997 8783 6055 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 19613 8823 19671 8829
rect 19613 8789 19625 8823
rect 19659 8820 19671 8823
rect 19978 8820 19984 8832
rect 19659 8792 19984 8820
rect 19659 8789 19671 8792
rect 19613 8783 19671 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8585 1823 8619
rect 1765 8579 1823 8585
rect 1780 8548 1808 8579
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 11146 8616 11152 8628
rect 2096 8588 11152 8616
rect 2096 8576 2102 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15804 8588 16037 8616
rect 15804 8576 15810 8588
rect 16025 8585 16037 8588
rect 16071 8616 16083 8619
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16071 8588 17049 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 2654 8551 2712 8557
rect 2654 8548 2666 8551
rect 1780 8520 2666 8548
rect 2654 8517 2666 8520
rect 2700 8517 2712 8551
rect 2654 8511 2712 8517
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 5776 8520 6469 8548
rect 5776 8508 5782 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 6914 8548 6920 8560
rect 6503 8520 6920 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7742 8548 7748 8560
rect 7703 8520 7748 8548
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 8110 8548 8116 8560
rect 8071 8520 8116 8548
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 11992 8548 12020 8576
rect 11716 8520 12020 8548
rect 11716 8492 11744 8520
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13326 8551 13384 8557
rect 13326 8548 13338 8551
rect 13228 8520 13338 8548
rect 13228 8508 13234 8520
rect 13326 8517 13338 8520
rect 13372 8517 13384 8551
rect 17052 8548 17080 8579
rect 19058 8576 19064 8628
rect 19116 8616 19122 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 19116 8588 19441 8616
rect 19116 8576 19122 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 18046 8548 18052 8560
rect 13326 8511 13384 8517
rect 15948 8520 16896 8548
rect 17052 8520 18052 8548
rect 15948 8492 15976 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2498 8480 2504 8492
rect 2455 8452 2504 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5960 8452 6377 8480
rect 5960 8440 5966 8452
rect 6365 8449 6377 8452
rect 6411 8480 6423 8483
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 6411 8452 7941 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7929 8449 7941 8452
rect 7975 8480 7987 8483
rect 8662 8480 8668 8492
rect 7975 8452 8668 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10226 8480 10232 8492
rect 10183 8452 10232 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 11698 8480 11704 8492
rect 11611 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 15841 8483 15899 8489
rect 12032 8452 12077 8480
rect 12032 8440 12038 8452
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 15930 8480 15936 8492
rect 15887 8452 15936 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16666 8480 16672 8492
rect 16627 8452 16672 8480
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16868 8489 16896 8520
rect 18046 8508 18052 8520
rect 18104 8548 18110 8560
rect 18782 8548 18788 8560
rect 18104 8520 18184 8548
rect 18104 8508 18110 8520
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17310 8480 17316 8492
rect 17175 8452 17316 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 18156 8489 18184 8520
rect 18432 8520 18788 8548
rect 18432 8489 18460 8520
rect 18782 8508 18788 8520
rect 18840 8548 18846 8560
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 18840 8520 19809 8548
rect 18840 8508 18846 8520
rect 19797 8517 19809 8520
rect 19843 8548 19855 8551
rect 19978 8548 19984 8560
rect 19843 8520 19984 8548
rect 19843 8517 19855 8520
rect 19797 8511 19855 8517
rect 19978 8508 19984 8520
rect 20036 8548 20042 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 20036 8520 20729 8548
rect 20036 8508 20042 8520
rect 20717 8517 20729 8520
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19484 8452 19625 8480
rect 19484 8440 19490 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20438 8480 20444 8492
rect 19935 8452 20444 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10502 8412 10508 8424
rect 10459 8384 10508 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 13081 8415 13139 8421
rect 13081 8412 13093 8415
rect 11480 8384 13093 8412
rect 11480 8372 11486 8384
rect 13081 8381 13093 8384
rect 13127 8381 13139 8415
rect 19628 8412 19656 8443
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 20548 8412 20576 8443
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 20864 8452 20909 8480
rect 20864 8440 20870 8452
rect 19628 8384 20576 8412
rect 13081 8375 13139 8381
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 20349 8347 20407 8353
rect 20349 8344 20361 8347
rect 16264 8316 20361 8344
rect 16264 8304 16270 8316
rect 20349 8313 20361 8316
rect 20395 8313 20407 8347
rect 20349 8307 20407 8313
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 8110 8276 8116 8288
rect 4672 8248 8116 8276
rect 4672 8236 4678 8248
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 13078 8276 13084 8288
rect 8352 8248 13084 8276
rect 8352 8236 8358 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 14458 8276 14464 8288
rect 14419 8248 14464 8276
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 2004 8044 2513 8072
rect 2004 8032 2010 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2501 8035 2559 8041
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4028 8044 7696 8072
rect 4028 8032 4034 8044
rect 7668 8004 7696 8044
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7800 8044 8125 8072
rect 7800 8032 7806 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10560 8044 10793 8072
rect 10560 8032 10566 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 11149 8075 11207 8081
rect 11149 8041 11161 8075
rect 11195 8072 11207 8075
rect 11882 8072 11888 8084
rect 11195 8044 11888 8072
rect 11195 8041 11207 8044
rect 11149 8035 11207 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12805 8075 12863 8081
rect 12805 8041 12817 8075
rect 12851 8072 12863 8075
rect 13354 8072 13360 8084
rect 12851 8044 13360 8072
rect 12851 8041 12863 8044
rect 12805 8035 12863 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 8294 8004 8300 8016
rect 7668 7976 8300 8004
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 13078 7964 13084 8016
rect 13136 8004 13142 8016
rect 13136 7976 13492 8004
rect 13136 7964 13142 7976
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3234 7936 3240 7948
rect 3191 7908 3240 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 8202 7896 8208 7948
rect 8260 7936 8266 7948
rect 8260 7908 11100 7936
rect 8260 7896 8266 7908
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1412 7800 1440 7831
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6604 7840 6745 7868
rect 6604 7828 6610 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10778 7868 10784 7880
rect 10376 7840 10784 7868
rect 10376 7828 10382 7840
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10962 7868 10968 7880
rect 10923 7840 10968 7868
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 7000 7803 7058 7809
rect 1412 7772 6960 7800
rect 1578 7732 1584 7744
rect 1539 7704 1584 7732
rect 1578 7692 1584 7704
rect 1636 7692 1642 7744
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3786 7732 3792 7744
rect 2915 7704 3792 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 6932 7732 6960 7772
rect 7000 7769 7012 7803
rect 7046 7800 7058 7803
rect 7098 7800 7104 7812
rect 7046 7772 7104 7800
rect 7046 7769 7058 7772
rect 7000 7763 7058 7769
rect 7098 7760 7104 7772
rect 7156 7760 7162 7812
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 11072 7800 11100 7908
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 13464 7945 13492 7976
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 11204 7908 13277 7936
rect 11204 7896 11210 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 16482 7936 16488 7948
rect 13495 7908 16488 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 17862 7936 17868 7948
rect 17823 7908 17868 7936
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 19978 7936 19984 7948
rect 19628 7908 19984 7936
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 17184 7840 17601 7868
rect 17184 7828 17190 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 17880 7868 17908 7896
rect 19426 7868 19432 7880
rect 17880 7840 19432 7868
rect 17589 7831 17647 7837
rect 19352 7834 19432 7840
rect 19426 7828 19432 7834
rect 19484 7828 19490 7880
rect 19628 7877 19656 7908
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 20530 7868 20536 7880
rect 19751 7840 20536 7868
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 19245 7803 19303 7809
rect 19245 7800 19257 7803
rect 8628 7772 10732 7800
rect 11072 7772 19257 7800
rect 8628 7760 8634 7772
rect 10594 7732 10600 7744
rect 6932 7704 10600 7732
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 10704 7732 10732 7772
rect 19245 7769 19257 7772
rect 19291 7769 19303 7803
rect 19245 7763 19303 7769
rect 13078 7732 13084 7744
rect 10704 7704 13084 7732
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 13814 7732 13820 7744
rect 13219 7704 13820 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 15010 7732 15016 7744
rect 14424 7704 15016 7732
rect 14424 7692 14430 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 3050 7528 3056 7540
rect 2179 7500 3056 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5902 7528 5908 7540
rect 5215 7500 5908 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 7984 7500 13461 7528
rect 7984 7488 7990 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13814 7528 13820 7540
rect 13449 7491 13507 7497
rect 13556 7500 13820 7528
rect 2593 7463 2651 7469
rect 2593 7429 2605 7463
rect 2639 7460 2651 7463
rect 2866 7460 2872 7472
rect 2639 7432 2872 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 4614 7460 4620 7472
rect 3252 7432 4620 7460
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2464 7364 2513 7392
rect 2464 7352 2470 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3252 7392 3280 7432
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 7466 7420 7472 7472
rect 7524 7460 7530 7472
rect 13081 7463 13139 7469
rect 7524 7432 12434 7460
rect 7524 7420 7530 7432
rect 2731 7364 3280 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 4045 7395 4103 7401
rect 4045 7392 4057 7395
rect 3384 7364 4057 7392
rect 3384 7352 3390 7364
rect 4045 7361 4057 7364
rect 4091 7361 4103 7395
rect 4045 7355 4103 7361
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6052 7364 6377 7392
rect 6052 7352 6058 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6549 7355 6607 7361
rect 1946 7324 1952 7336
rect 1907 7296 1952 7324
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 3200 7296 3801 7324
rect 3200 7284 3206 7296
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3804 7188 3832 7287
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 6564 7324 6592 7355
rect 6914 7352 6920 7364
rect 6972 7392 6978 7404
rect 7282 7392 7288 7404
rect 6972 7364 7288 7392
rect 6972 7352 6978 7364
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 7892 7364 8585 7392
rect 7892 7352 7898 7364
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 8846 7392 8852 7404
rect 8720 7364 8765 7392
rect 8807 7364 8852 7392
rect 8720 7352 8726 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 4856 7296 6592 7324
rect 6641 7327 6699 7333
rect 4856 7284 4862 7296
rect 6641 7293 6653 7327
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 9766 7324 9772 7336
rect 6779 7296 9772 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 6656 7256 6684 7287
rect 9766 7284 9772 7296
rect 9824 7324 9830 7336
rect 10520 7324 10548 7355
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10652 7364 10697 7392
rect 10652 7352 10658 7364
rect 10778 7324 10784 7336
rect 9824 7296 10784 7324
rect 9824 7284 9830 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 12406 7324 12434 7432
rect 13081 7429 13093 7463
rect 13127 7460 13139 7463
rect 13556 7460 13584 7500
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 14458 7528 14464 7540
rect 13872 7500 14464 7528
rect 13872 7488 13878 7500
rect 14458 7488 14464 7500
rect 14516 7528 14522 7540
rect 14921 7531 14979 7537
rect 14921 7528 14933 7531
rect 14516 7500 14933 7528
rect 14516 7488 14522 7500
rect 14921 7497 14933 7500
rect 14967 7497 14979 7531
rect 18782 7528 18788 7540
rect 18743 7500 18788 7528
rect 14921 7491 14979 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 13127 7432 13584 7460
rect 13832 7432 17448 7460
rect 13127 7429 13139 7432
rect 13081 7423 13139 7429
rect 13832 7404 13860 7432
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 13170 7392 13176 7404
rect 13131 7364 13176 7392
rect 12897 7355 12955 7361
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12406 7296 12725 7324
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 5500 7228 6684 7256
rect 9217 7259 9275 7265
rect 5500 7216 5506 7228
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 12912 7256 12940 7355
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13814 7392 13820 7404
rect 13679 7364 13820 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7392 13967 7395
rect 14642 7392 14648 7404
rect 13955 7364 14648 7392
rect 13955 7361 13967 7364
rect 13909 7355 13967 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 14752 7401 14780 7432
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 14737 7355 14795 7361
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 17420 7401 17448 7432
rect 17405 7395 17463 7401
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17451 7364 18613 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19242 7392 19248 7404
rect 18923 7364 19248 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 13078 7284 13084 7336
rect 13136 7324 13142 7336
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 13136 7296 14565 7324
rect 13136 7284 13142 7296
rect 14553 7293 14565 7296
rect 14599 7293 14611 7327
rect 17126 7324 17132 7336
rect 17087 7296 17132 7324
rect 14553 7287 14611 7293
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 13814 7256 13820 7268
rect 9263 7228 12434 7256
rect 12912 7228 13820 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 6546 7188 6552 7200
rect 3804 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10870 7188 10876 7200
rect 10831 7160 10876 7188
rect 10870 7148 10876 7160
rect 10928 7148 10934 7200
rect 12406 7188 12434 7228
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14200 7228 14504 7256
rect 14200 7188 14228 7228
rect 12406 7160 14228 7188
rect 14277 7191 14335 7197
rect 14277 7157 14289 7191
rect 14323 7188 14335 7191
rect 14366 7188 14372 7200
rect 14323 7160 14372 7188
rect 14323 7157 14335 7160
rect 14277 7151 14335 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14476 7188 14504 7228
rect 15746 7188 15752 7200
rect 14476 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 18414 7188 18420 7200
rect 18375 7160 18420 7188
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 2866 6984 2872 6996
rect 2779 6956 2872 6984
rect 2866 6944 2872 6956
rect 2924 6984 2930 6996
rect 4062 6984 4068 6996
rect 2924 6956 4068 6984
rect 2924 6944 2930 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 6052 6956 6101 6984
rect 6052 6944 6058 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7834 6984 7840 6996
rect 7423 6956 7840 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 7944 6956 12434 6984
rect 7285 6919 7343 6925
rect 7285 6916 7297 6919
rect 7116 6888 7297 6916
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 2004 6820 6040 6848
rect 2004 6808 2010 6820
rect 6012 6792 6040 6820
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7116 6848 7144 6888
rect 7285 6885 7297 6888
rect 7331 6885 7343 6919
rect 7285 6879 7343 6885
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 7944 6916 7972 6956
rect 7708 6888 7972 6916
rect 12406 6916 12434 6956
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13228 6956 22094 6984
rect 13228 6944 13234 6956
rect 18414 6916 18420 6928
rect 12406 6888 18420 6916
rect 7708 6876 7714 6888
rect 18414 6876 18420 6888
rect 18472 6876 18478 6928
rect 22066 6916 22094 6956
rect 37274 6916 37280 6928
rect 22066 6888 37280 6916
rect 37274 6876 37280 6888
rect 37332 6876 37338 6928
rect 6788 6820 7144 6848
rect 7193 6851 7251 6857
rect 6788 6808 6794 6820
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 8846 6848 8852 6860
rect 7239 6820 8852 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 14277 6851 14335 6857
rect 9232 6820 9536 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 3970 6780 3976 6792
rect 1719 6752 3976 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4614 6780 4620 6792
rect 4571 6752 4620 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5442 6780 5448 6792
rect 4847 6752 5448 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5994 6780 6000 6792
rect 5907 6752 6000 6780
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6104 6752 7113 6780
rect 2406 6672 2412 6724
rect 2464 6712 2470 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2464 6684 2697 6712
rect 2464 6672 2470 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 3510 6672 3516 6724
rect 3568 6712 3574 6724
rect 6104 6712 6132 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 3568 6684 6132 6712
rect 3568 6672 3574 6684
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 2885 6647 2943 6653
rect 2885 6644 2897 6647
rect 2832 6616 2897 6644
rect 2832 6604 2838 6616
rect 2885 6613 2897 6616
rect 2931 6613 2943 6647
rect 2885 6607 2943 6613
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 4798 6644 4804 6656
rect 3099 6616 4804 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7116 6644 7144 6743
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7340 6752 7573 6780
rect 7340 6740 7346 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 9232 6780 9260 6820
rect 9508 6789 9536 6820
rect 14277 6817 14289 6851
rect 14323 6848 14335 6851
rect 14458 6848 14464 6860
rect 14323 6820 14464 6848
rect 14323 6817 14335 6820
rect 14277 6811 14335 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 15804 6820 15853 6848
rect 15804 6808 15810 6820
rect 15841 6817 15853 6820
rect 15887 6848 15899 6851
rect 17126 6848 17132 6860
rect 15887 6820 17132 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 7708 6752 9260 6780
rect 9309 6783 9367 6789
rect 7708 6740 7714 6752
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 9493 6743 9551 6749
rect 9324 6712 9352 6743
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 14550 6780 14556 6792
rect 14511 6752 14556 6780
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 15988 6752 16129 6780
rect 15988 6740 15994 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 10312 6715 10370 6721
rect 9324 6684 9536 6712
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 7116 6616 9413 6644
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9508 6644 9536 6684
rect 10312 6681 10324 6715
rect 10358 6712 10370 6715
rect 10410 6712 10416 6724
rect 10358 6684 10416 6712
rect 10358 6681 10370 6684
rect 10312 6675 10370 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 16132 6712 16160 6743
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 17405 6783 17463 6789
rect 17405 6780 17417 6783
rect 16264 6752 17417 6780
rect 16264 6740 16270 6752
rect 17405 6749 17417 6752
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 16298 6712 16304 6724
rect 16132 6684 16304 6712
rect 16298 6672 16304 6684
rect 16356 6672 16362 6724
rect 10502 6644 10508 6656
rect 9508 6616 10508 6644
rect 9401 6607 9459 6613
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10652 6616 11437 6644
rect 10652 6604 10658 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 3697 6443 3755 6449
rect 3697 6440 3709 6443
rect 2823 6412 3709 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 3697 6409 3709 6412
rect 3743 6409 3755 6443
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 3697 6403 3755 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10781 6443 10839 6449
rect 10781 6409 10793 6443
rect 10827 6440 10839 6443
rect 10870 6440 10876 6452
rect 10827 6412 10876 6440
rect 10827 6409 10839 6412
rect 10781 6403 10839 6409
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 14550 6440 14556 6452
rect 14507 6412 14556 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 14550 6400 14556 6412
rect 14608 6440 14614 6452
rect 15286 6440 15292 6452
rect 14608 6412 15292 6440
rect 14608 6400 14614 6412
rect 15286 6400 15292 6412
rect 15344 6440 15350 6452
rect 15381 6443 15439 6449
rect 15381 6440 15393 6443
rect 15344 6412 15393 6440
rect 15344 6400 15350 6412
rect 15381 6409 15393 6412
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6409 16911 6443
rect 16853 6403 16911 6409
rect 3326 6372 3332 6384
rect 3287 6344 3332 6372
rect 3326 6332 3332 6344
rect 3384 6332 3390 6384
rect 5994 6332 6000 6384
rect 6052 6372 6058 6384
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6052 6344 7113 6372
rect 6052 6332 6058 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7285 6375 7343 6381
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 7374 6372 7380 6384
rect 7331 6344 7380 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 7374 6332 7380 6344
rect 7432 6332 7438 6384
rect 11330 6372 11336 6384
rect 10612 6344 11336 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 2774 6304 2780 6316
rect 2731 6276 2780 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 1412 6168 1440 6267
rect 2700 6168 2728 6267
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 3510 6304 3516 6316
rect 3471 6276 3516 6304
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 10612 6313 10640 6344
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 11698 6372 11704 6384
rect 11388 6344 11704 6372
rect 11388 6332 11394 6344
rect 11698 6332 11704 6344
rect 11756 6332 11762 6384
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 13504 6344 15025 6372
rect 13504 6332 13510 6344
rect 15013 6341 15025 6344
rect 15059 6341 15071 6375
rect 15654 6372 15660 6384
rect 15013 6335 15071 6341
rect 15212 6344 15660 6372
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6273 10655 6307
rect 10870 6304 10876 6316
rect 10831 6276 10876 6304
rect 10597 6267 10655 6273
rect 3234 6196 3240 6248
rect 3292 6236 3298 6248
rect 3804 6236 3832 6267
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 15212 6313 15240 6344
rect 15654 6332 15660 6344
rect 15712 6372 15718 6384
rect 16206 6372 16212 6384
rect 15712 6344 16212 6372
rect 15712 6332 15718 6344
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16868 6372 16896 6403
rect 17742 6375 17800 6381
rect 17742 6372 17754 6375
rect 16868 6344 17754 6372
rect 17742 6341 17754 6344
rect 17788 6341 17800 6375
rect 17742 6335 17800 6341
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13872 6276 14289 6304
rect 13872 6264 13878 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6273 15255 6307
rect 15197 6267 15255 6273
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 16022 6304 16028 6316
rect 15519 6276 16028 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 3292 6208 3832 6236
rect 3292 6196 3298 6208
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 7248 6208 14105 6236
rect 7248 6196 7254 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14568 6236 14596 6267
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16448 6276 17049 6304
rect 16448 6264 16454 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 38562 6304 38568 6316
rect 17037 6267 17095 6273
rect 17420 6276 38568 6304
rect 17420 6236 17448 6276
rect 38562 6264 38568 6276
rect 38620 6264 38626 6316
rect 14568 6208 17448 6236
rect 17497 6239 17555 6245
rect 14093 6199 14151 6205
rect 17497 6205 17509 6239
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 5258 6168 5264 6180
rect 1412 6140 2636 6168
rect 2700 6140 5264 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2608 6100 2636 6140
rect 5258 6128 5264 6140
rect 5316 6128 5322 6180
rect 10686 6168 10692 6180
rect 7116 6140 10692 6168
rect 7116 6100 7144 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 16850 6128 16856 6180
rect 16908 6168 16914 6180
rect 17512 6168 17540 6199
rect 16908 6140 17540 6168
rect 16908 6128 16914 6140
rect 18874 6100 18880 6112
rect 2608 6072 7144 6100
rect 18835 6072 18880 6100
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4028 5868 7512 5896
rect 4028 5856 4034 5868
rect 7484 5828 7512 5868
rect 9950 5856 9956 5908
rect 10008 5896 10014 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 10008 5868 14473 5896
rect 10008 5856 10014 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15252 5868 15485 5896
rect 15252 5856 15258 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 15473 5859 15531 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 7484 5800 12434 5828
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3234 5760 3240 5772
rect 3099 5732 3240 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 6546 5760 6552 5772
rect 6507 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 12406 5760 12434 5800
rect 16482 5788 16488 5840
rect 16540 5828 16546 5840
rect 16540 5800 16988 5828
rect 16540 5788 16546 5800
rect 16960 5769 16988 5800
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 12406 5732 16865 5760
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16853 5723 16911 5729
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 6822 5701 6828 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 1728 5664 3801 5692
rect 1728 5652 1734 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 6816 5692 6828 5701
rect 6783 5664 6828 5692
rect 3789 5655 3847 5661
rect 6816 5655 6828 5664
rect 6822 5652 6828 5655
rect 6880 5652 6886 5704
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5692 14979 5695
rect 15010 5692 15016 5704
rect 14967 5664 15016 5692
rect 14967 5661 14979 5664
rect 14921 5655 14979 5661
rect 2869 5627 2927 5633
rect 2869 5624 2881 5627
rect 1412 5596 2881 5624
rect 1412 5565 1440 5596
rect 2869 5593 2881 5596
rect 2915 5593 2927 5627
rect 2869 5587 2927 5593
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5525 1455 5559
rect 1397 5519 1455 5525
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2590 5556 2596 5568
rect 2455 5528 2596 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 3602 5556 3608 5568
rect 2823 5528 3608 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 6730 5556 6736 5568
rect 6236 5528 6736 5556
rect 6236 5516 6242 5528
rect 6730 5516 6736 5528
rect 6788 5556 6794 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 6788 5528 7941 5556
rect 6788 5516 6794 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 14660 5556 14688 5655
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15378 5652 15384 5704
rect 15436 5692 15442 5704
rect 15654 5692 15660 5704
rect 15436 5664 15660 5692
rect 15436 5652 15442 5664
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15930 5692 15936 5704
rect 15891 5664 15936 5692
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 14829 5627 14887 5633
rect 14829 5593 14841 5627
rect 14875 5624 14887 5627
rect 15286 5624 15292 5636
rect 14875 5596 15292 5624
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15378 5556 15384 5568
rect 14660 5528 15384 5556
rect 7929 5519 7987 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16758 5556 16764 5568
rect 15887 5528 16764 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5321 1455 5355
rect 3602 5352 3608 5364
rect 3563 5324 3608 5352
rect 1397 5315 1455 5321
rect 1412 5284 1440 5315
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 10744 5324 12909 5352
rect 10744 5312 10750 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 13596 5324 14289 5352
rect 13596 5312 13602 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 15160 5324 15209 5352
rect 15160 5312 15166 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 15197 5315 15255 5321
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 15896 5324 16681 5352
rect 15896 5312 15902 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 17770 5312 17776 5364
rect 17828 5352 17834 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 17828 5324 18613 5352
rect 17828 5312 17834 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 18601 5315 18659 5321
rect 6822 5284 6828 5296
rect 1412 5256 6828 5284
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 14645 5287 14703 5293
rect 14645 5253 14657 5287
rect 14691 5284 14703 5287
rect 15286 5284 15292 5296
rect 14691 5256 15292 5284
rect 14691 5253 14703 5256
rect 14645 5247 14703 5253
rect 15286 5244 15292 5256
rect 15344 5284 15350 5296
rect 15565 5287 15623 5293
rect 15565 5284 15577 5287
rect 15344 5256 15577 5284
rect 15344 5244 15350 5256
rect 15565 5253 15577 5256
rect 15611 5253 15623 5287
rect 15565 5247 15623 5253
rect 16758 5244 16764 5296
rect 16816 5284 16822 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 16816 5256 17049 5284
rect 16816 5244 16822 5256
rect 17037 5253 17049 5256
rect 17083 5284 17095 5287
rect 18874 5284 18880 5296
rect 17083 5256 18880 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 18969 5287 19027 5293
rect 18969 5253 18981 5287
rect 19015 5284 19027 5287
rect 19334 5284 19340 5296
rect 19015 5256 19340 5284
rect 19015 5253 19027 5256
rect 18969 5247 19027 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2314 5216 2320 5228
rect 2271 5188 2320 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2498 5225 2504 5228
rect 2492 5179 2504 5225
rect 2556 5216 2562 5228
rect 4249 5219 4307 5225
rect 2556 5188 2592 5216
rect 2498 5176 2504 5179
rect 2556 5176 2562 5188
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4614 5216 4620 5228
rect 4295 5188 4620 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5442 5216 5448 5228
rect 4939 5188 5448 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5442 5176 5448 5188
rect 5500 5216 5506 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5500 5188 6561 5216
rect 5500 5176 5506 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 6549 5179 6607 5185
rect 9766 5176 9772 5188
rect 9824 5216 9830 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 9824 5188 10609 5216
rect 9824 5176 9830 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10744 5188 10789 5216
rect 10744 5176 10750 5188
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11773 5219 11831 5225
rect 11773 5216 11785 5219
rect 11204 5188 11785 5216
rect 11204 5176 11210 5188
rect 11773 5185 11785 5188
rect 11819 5185 11831 5219
rect 11773 5179 11831 5185
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14737 5219 14795 5225
rect 14737 5185 14749 5219
rect 14783 5216 14795 5219
rect 15102 5216 15108 5228
rect 14783 5188 15108 5216
rect 14783 5185 14795 5188
rect 14737 5179 14795 5185
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 3844 5120 4721 5148
rect 3844 5108 3850 5120
rect 4709 5117 4721 5120
rect 4755 5117 4767 5151
rect 4709 5111 4767 5117
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5117 6423 5151
rect 9858 5148 9864 5160
rect 9819 5120 9864 5148
rect 6365 5111 6423 5117
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 6380 5080 6408 5111
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 10100 5120 11529 5148
rect 10100 5108 10106 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 14476 5148 14504 5179
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 15378 5216 15384 5228
rect 15339 5188 15384 5216
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 15654 5176 15660 5228
rect 15712 5216 15718 5228
rect 16850 5216 16856 5228
rect 15712 5188 15757 5216
rect 16811 5188 16856 5216
rect 15712 5176 15718 5188
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 18782 5216 18788 5228
rect 18743 5188 18788 5216
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 19061 5219 19119 5225
rect 19061 5185 19073 5219
rect 19107 5216 19119 5219
rect 30282 5216 30288 5228
rect 19107 5188 30288 5216
rect 19107 5185 19119 5188
rect 19061 5179 19119 5185
rect 30282 5176 30288 5188
rect 30340 5176 30346 5228
rect 15396 5148 15424 5176
rect 14476 5120 15424 5148
rect 11517 5111 11575 5117
rect 10502 5080 10508 5092
rect 3936 5052 6408 5080
rect 9968 5052 10508 5080
rect 3936 5040 3942 5052
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5718 5012 5724 5024
rect 5123 4984 5724 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 8202 5012 8208 5024
rect 6779 4984 8208 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9968 5021 9996 5052
rect 10502 5040 10508 5052
rect 10560 5080 10566 5092
rect 10560 5052 10640 5080
rect 10560 5040 10566 5052
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 4981 10011 5015
rect 10134 5012 10140 5024
rect 10095 4984 10140 5012
rect 9953 4975 10011 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10612 5021 10640 5052
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11514 5012 11520 5024
rect 11011 4984 11520 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2498 4808 2504 4820
rect 2455 4780 2504 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 9858 4808 9864 4820
rect 2746 4780 9864 4808
rect 2746 4740 2774 4780
rect 9858 4768 9864 4780
rect 9916 4808 9922 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 9916 4780 10333 4808
rect 9916 4768 9922 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 11146 4808 11152 4820
rect 11107 4780 11152 4808
rect 10321 4771 10379 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15381 4811 15439 4817
rect 15381 4808 15393 4811
rect 14884 4780 15393 4808
rect 14884 4768 14890 4780
rect 15381 4777 15393 4780
rect 15427 4777 15439 4811
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 15381 4771 15439 4777
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 1412 4712 2774 4740
rect 1412 4613 1440 4712
rect 5442 4700 5448 4752
rect 5500 4700 5506 4752
rect 3602 4632 3608 4684
rect 3660 4672 3666 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3660 4644 3801 4672
rect 3660 4632 3666 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 5460 4672 5488 4700
rect 3789 4635 3847 4641
rect 3988 4644 6316 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 1397 4567 1455 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3988 4613 4016 4644
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3200 4576 3249 4604
rect 3200 4564 3206 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 4212 4576 4629 4604
rect 4212 4564 4218 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 6288 4613 6316 4644
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 6604 4644 8953 4672
rect 6604 4632 6610 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 16577 4675 16635 4681
rect 16577 4672 16589 4675
rect 8941 4635 8999 4641
rect 15580 4644 16589 4672
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 5224 4576 5457 4604
rect 5224 4564 5230 4576
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 8956 4604 8984 4635
rect 10042 4604 10048 4616
rect 8956 4576 10048 4604
rect 6273 4567 6331 4573
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 6104 4536 6132 4567
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 11330 4604 11336 4616
rect 11291 4576 11336 4604
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11514 4604 11520 4616
rect 11475 4576 11520 4604
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 15580 4613 15608 4644
rect 16577 4641 16589 4644
rect 16623 4672 16635 4675
rect 16850 4672 16856 4684
rect 16623 4644 16856 4672
rect 16623 4641 16635 4644
rect 16577 4635 16635 4641
rect 16850 4632 16856 4644
rect 16908 4672 16914 4684
rect 18782 4672 18788 4684
rect 16908 4644 18788 4672
rect 16908 4632 16914 4644
rect 15565 4607 15623 4613
rect 11664 4576 11709 4604
rect 11664 4564 11670 4576
rect 15565 4573 15577 4607
rect 15611 4573 15623 4607
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15565 4567 15623 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 16298 4604 16304 4616
rect 16259 4576 16304 4604
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 18432 4613 18460 4644
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 18932 4644 19257 4672
rect 18932 4632 18938 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 19058 4604 19064 4616
rect 18739 4576 19064 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 19521 4567 19579 4573
rect 5408 4508 6132 4536
rect 9208 4539 9266 4545
rect 5408 4496 5414 4508
rect 9208 4505 9220 4539
rect 9254 4536 9266 4539
rect 9766 4536 9772 4548
rect 9254 4508 9772 4536
rect 9254 4505 9266 4508
rect 9208 4499 9266 4505
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 15749 4539 15807 4545
rect 15749 4505 15761 4539
rect 15795 4536 15807 4539
rect 16758 4536 16764 4548
rect 15795 4508 16764 4536
rect 15795 4505 15807 4508
rect 15749 4499 15807 4505
rect 16758 4496 16764 4508
rect 16816 4496 16822 4548
rect 19334 4536 19340 4548
rect 18616 4508 19340 4536
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4157 4471 4215 4477
rect 4157 4437 4169 4471
rect 4203 4468 4215 4471
rect 4338 4468 4344 4480
rect 4203 4440 4344 4468
rect 4203 4437 4215 4440
rect 4157 4431 4215 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 10226 4468 10232 4480
rect 6503 4440 10232 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 18506 4428 18512 4480
rect 18564 4468 18570 4480
rect 18616 4477 18644 4508
rect 19334 4496 19340 4508
rect 19392 4536 19398 4548
rect 19536 4536 19564 4567
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 19392 4508 19564 4536
rect 19392 4496 19398 4508
rect 18601 4471 18659 4477
rect 18601 4468 18613 4471
rect 18564 4440 18613 4468
rect 18564 4428 18570 4440
rect 18601 4437 18613 4440
rect 18647 4437 18659 4471
rect 18601 4431 18659 4437
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4468 24455 4471
rect 24670 4468 24676 4480
rect 24443 4440 24676 4468
rect 24443 4437 24455 4440
rect 24397 4431 24455 4437
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10226 4224 10232 4276
rect 10284 4264 10290 4276
rect 24578 4264 24584 4276
rect 10284 4236 24584 4264
rect 10284 4224 10290 4236
rect 24578 4224 24584 4236
rect 24636 4224 24642 4276
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7926 4196 7932 4208
rect 6779 4168 7932 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 18506 4156 18512 4208
rect 18564 4196 18570 4208
rect 18969 4199 19027 4205
rect 18969 4196 18981 4199
rect 18564 4168 18981 4196
rect 18564 4156 18570 4168
rect 18969 4165 18981 4168
rect 19015 4196 19027 4199
rect 19889 4199 19947 4205
rect 19889 4196 19901 4199
rect 19015 4168 19901 4196
rect 19015 4165 19027 4168
rect 18969 4159 19027 4165
rect 19889 4165 19901 4168
rect 19935 4165 19947 4199
rect 19889 4159 19947 4165
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1443 4100 2268 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 2240 4001 2268 4100
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 2372 4100 2421 4128
rect 2372 4088 2378 4100
rect 2409 4097 2421 4100
rect 2455 4128 2467 4131
rect 3142 4128 3148 4140
rect 2455 4100 3148 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3292 4100 3433 4128
rect 3292 4088 3298 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 3620 4060 3648 4091
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 4338 4128 4344 4140
rect 3752 4100 3797 4128
rect 4299 4100 4344 4128
rect 3752 4088 3758 4100
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 2740 4032 3648 4060
rect 2740 4020 2746 4032
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 5644 4060 5672 4091
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 9766 4128 9772 4140
rect 6880 4100 6925 4128
rect 9727 4100 9772 4128
rect 6880 4088 6886 4100
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 9953 4091 10011 4097
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 4028 4032 5672 4060
rect 5736 4032 6929 4060
rect 4028 4020 4034 4032
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3961 2283 3995
rect 2225 3955 2283 3961
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 3660 3964 4997 3992
rect 3660 3952 3666 3964
rect 4985 3961 4997 3964
rect 5031 3961 5043 3995
rect 4985 3955 5043 3961
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 5445 3995 5503 4001
rect 5445 3992 5457 3995
rect 5316 3964 5457 3992
rect 5316 3952 5322 3964
rect 5445 3961 5457 3964
rect 5491 3961 5503 3995
rect 5445 3955 5503 3961
rect 198 3884 204 3936
rect 256 3924 262 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 256 3896 1593 3924
rect 256 3884 262 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3878 3924 3884 3936
rect 3283 3896 3884 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4706 3924 4712 3936
rect 4203 3896 4712 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5074 3884 5080 3936
rect 5132 3924 5138 3936
rect 5736 3924 5764 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 9968 4060 9996 4091
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 11296 4100 14289 4128
rect 11296 4088 11302 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 14277 4091 14335 4097
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 18782 4128 18788 4140
rect 18743 4100 18788 4128
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 11330 4060 11336 4072
rect 9968 4032 11336 4060
rect 6917 4023 6975 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 16298 4020 16304 4072
rect 16356 4060 16362 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 16356 4032 16681 4060
rect 16356 4020 16362 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 16945 4063 17003 4069
rect 16945 4029 16957 4063
rect 16991 4060 17003 4063
rect 17586 4060 17592 4072
rect 16991 4032 17592 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 19076 4060 19104 4091
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19484 4100 19533 4128
rect 19484 4088 19490 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19702 4128 19708 4140
rect 19663 4100 19708 4128
rect 19521 4091 19579 4097
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4128 20039 4131
rect 25590 4128 25596 4140
rect 20027 4100 25596 4128
rect 20027 4097 20039 4100
rect 19981 4091 20039 4097
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 28810 4060 28816 4072
rect 19076 4032 28816 4060
rect 28810 4020 28816 4032
rect 28868 4020 28874 4072
rect 10962 3952 10968 4004
rect 11020 3992 11026 4004
rect 21266 3992 21272 4004
rect 11020 3964 21272 3992
rect 11020 3952 11026 3964
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 5132 3896 5764 3924
rect 6365 3927 6423 3933
rect 5132 3884 5138 3896
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6454 3924 6460 3936
rect 6411 3896 6460 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 11882 3924 11888 3936
rect 8444 3896 11888 3924
rect 8444 3884 8450 3896
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14826 3924 14832 3936
rect 14139 3896 14832 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 4798 3720 4804 3732
rect 2746 3692 4804 3720
rect 658 3612 664 3664
rect 716 3652 722 3664
rect 2593 3655 2651 3661
rect 2593 3652 2605 3655
rect 716 3624 2605 3652
rect 716 3612 722 3624
rect 2593 3621 2605 3624
rect 2639 3621 2651 3655
rect 2593 3615 2651 3621
rect 2746 3584 2774 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11241 3723 11299 3729
rect 9640 3692 11100 3720
rect 9640 3680 9646 3692
rect 11072 3652 11100 3692
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 11606 3720 11612 3732
rect 11287 3692 11612 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 16574 3720 16580 3732
rect 16535 3692 16580 3720
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 18233 3723 18291 3729
rect 18233 3720 18245 3723
rect 17552 3692 18245 3720
rect 17552 3680 17558 3692
rect 18233 3689 18245 3692
rect 18279 3689 18291 3723
rect 18233 3683 18291 3689
rect 15746 3652 15752 3664
rect 11072 3624 15752 3652
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 57977 3655 58035 3661
rect 57977 3652 57989 3655
rect 16172 3624 57989 3652
rect 16172 3612 16178 3624
rect 57977 3621 57989 3624
rect 58023 3621 58035 3655
rect 57977 3615 58035 3621
rect 1688 3556 2774 3584
rect 1688 3525 1716 3556
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3200 3556 3801 3584
rect 3200 3544 3206 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 10778 3544 10784 3596
rect 10836 3584 10842 3596
rect 14645 3587 14703 3593
rect 10836 3556 11836 3584
rect 10836 3544 10842 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 3050 3516 3056 3528
rect 2455 3488 3056 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4045 3519 4103 3525
rect 4045 3516 4057 3519
rect 3936 3488 4057 3516
rect 3936 3476 3942 3488
rect 4045 3485 4057 3488
rect 4091 3485 4103 3519
rect 4045 3479 4103 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3485 5871 3519
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 5813 3479 5871 3485
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 5828 3448 5856 3479
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7524 3488 7757 3516
rect 7524 3476 7530 3488
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10468 3488 10701 3516
rect 10468 3476 10474 3488
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 11422 3516 11428 3528
rect 11383 3488 11428 3516
rect 10689 3479 10747 3485
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 11624 3525 11652 3556
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11716 3448 11744 3479
rect 3752 3420 5856 3448
rect 7576 3420 11744 3448
rect 3752 3408 3758 3420
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1636 3352 1869 3380
rect 1636 3340 1642 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 1857 3343 1915 3349
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 5169 3383 5227 3389
rect 5169 3380 5181 3383
rect 2740 3352 5181 3380
rect 2740 3340 2746 3352
rect 5169 3349 5181 3352
rect 5215 3349 5227 3383
rect 6270 3380 6276 3392
rect 6231 3352 6276 3380
rect 5169 3343 5227 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 7576 3389 7604 3420
rect 6917 3383 6975 3389
rect 6917 3380 6929 3383
rect 6420 3352 6929 3380
rect 6420 3340 6426 3352
rect 6917 3349 6929 3352
rect 6963 3349 6975 3383
rect 6917 3343 6975 3349
rect 7561 3383 7619 3389
rect 7561 3349 7573 3383
rect 7607 3349 7619 3383
rect 7561 3343 7619 3349
rect 10505 3383 10563 3389
rect 10505 3349 10517 3383
rect 10551 3380 10563 3383
rect 10962 3380 10968 3392
rect 10551 3352 10968 3380
rect 10551 3349 10563 3352
rect 10505 3343 10563 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11808 3380 11836 3556
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 16298 3584 16304 3596
rect 14691 3556 16304 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 16942 3584 16948 3596
rect 16776 3556 16948 3584
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 12400 3488 12633 3516
rect 12400 3476 12406 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13412 3488 13553 3516
rect 13412 3476 13418 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14792 3488 14933 3516
rect 14792 3476 14798 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16206 3516 16212 3528
rect 16163 3488 16212 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16776 3525 16804 3556
rect 16942 3544 16948 3556
rect 17000 3584 17006 3596
rect 17586 3584 17592 3596
rect 17000 3556 17592 3584
rect 17000 3544 17006 3556
rect 17586 3544 17592 3556
rect 17644 3584 17650 3596
rect 19702 3584 19708 3596
rect 17644 3556 19708 3584
rect 17644 3544 17650 3556
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17037 3519 17095 3525
rect 17037 3485 17049 3519
rect 17083 3516 17095 3519
rect 18322 3516 18328 3528
rect 17083 3488 18328 3516
rect 17083 3485 17095 3488
rect 17037 3479 17095 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18432 3525 18460 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18564 3488 18613 3516
rect 18564 3476 18570 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 25682 3516 25688 3528
rect 18739 3488 25688 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 11882 3408 11888 3460
rect 11940 3448 11946 3460
rect 15194 3448 15200 3460
rect 11940 3420 15200 3448
rect 11940 3408 11946 3420
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 57793 3451 57851 3457
rect 57793 3417 57805 3451
rect 57839 3448 57851 3451
rect 59630 3448 59636 3460
rect 57839 3420 59636 3448
rect 57839 3417 57851 3420
rect 57793 3411 57851 3417
rect 59630 3408 59636 3420
rect 59688 3408 59694 3460
rect 12618 3380 12624 3392
rect 11808 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12768 3352 13369 3380
rect 12768 3340 12774 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 15933 3383 15991 3389
rect 15933 3380 15945 3383
rect 14976 3352 15945 3380
rect 14976 3340 14982 3352
rect 15933 3349 15945 3352
rect 15979 3349 15991 3383
rect 15933 3343 15991 3349
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 16945 3383 17003 3389
rect 16945 3380 16957 3383
rect 16724 3352 16957 3380
rect 16724 3340 16730 3352
rect 16945 3349 16957 3352
rect 16991 3380 17003 3383
rect 17034 3380 17040 3392
rect 16991 3352 17040 3380
rect 16991 3349 17003 3352
rect 16945 3343 17003 3349
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 19978 3380 19984 3392
rect 17184 3352 19984 3380
rect 17184 3340 17190 3352
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 4062 3176 4068 3188
rect 2188 3148 4068 3176
rect 2188 3136 2194 3148
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 7926 3176 7932 3188
rect 7839 3148 7932 3176
rect 7926 3136 7932 3148
rect 7984 3176 7990 3188
rect 10505 3179 10563 3185
rect 7984 3148 9067 3176
rect 7984 3136 7990 3148
rect 6178 3108 6184 3120
rect 3436 3080 6184 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1946 3040 1952 3052
rect 1719 3012 1952 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2682 3040 2688 3052
rect 2643 3012 2688 3040
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3436 3049 3464 3080
rect 6178 3068 6184 3080
rect 6236 3068 6242 3120
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 6794 3111 6852 3117
rect 6794 3108 6806 3111
rect 6328 3080 6806 3108
rect 6328 3068 6334 3080
rect 6794 3077 6806 3080
rect 6840 3077 6852 3111
rect 6794 3071 6852 3077
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4614 3040 4620 3052
rect 4479 3012 4620 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5718 3040 5724 3052
rect 4816 3012 5212 3040
rect 5679 3012 5724 3040
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 4816 2972 4844 3012
rect 2464 2944 4844 2972
rect 4893 2975 4951 2981
rect 2464 2932 2470 2944
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 5074 2972 5080 2984
rect 4939 2944 5080 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5184 2972 5212 3012
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8260 3012 8585 3040
rect 8260 3000 8266 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 6362 2972 6368 2984
rect 5184 2944 6368 2972
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 9039 2972 9067 3148
rect 10505 3145 10517 3179
rect 10551 3176 10563 3179
rect 10870 3176 10876 3188
rect 10551 3148 10876 3176
rect 10551 3145 10563 3148
rect 10505 3139 10563 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12032 3148 12265 3176
rect 12032 3136 12038 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 13998 3136 14004 3188
rect 14056 3176 14062 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14056 3148 14473 3176
rect 14056 3136 14062 3148
rect 14461 3145 14473 3148
rect 14507 3145 14519 3179
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 14461 3139 14519 3145
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 23661 3179 23719 3185
rect 23661 3176 23673 3179
rect 18380 3148 23673 3176
rect 18380 3136 18386 3148
rect 23661 3145 23673 3148
rect 23707 3145 23719 3179
rect 56965 3179 57023 3185
rect 56965 3176 56977 3179
rect 23661 3139 23719 3145
rect 26206 3148 56977 3176
rect 12618 3108 12624 3120
rect 10704 3080 11468 3108
rect 12531 3080 12624 3108
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9364 3012 10057 3040
rect 9364 3000 9370 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10704 3049 10732 3080
rect 11440 3052 11468 3080
rect 12618 3068 12624 3080
rect 12676 3108 12682 3120
rect 14829 3111 14887 3117
rect 14829 3108 14841 3111
rect 12676 3080 14841 3108
rect 12676 3068 12682 3080
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10652 3012 10701 3040
rect 10652 3000 10658 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10836 3012 10885 3040
rect 10836 3000 10842 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11020 3012 11065 3040
rect 11020 3000 11026 3012
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 12456 3043 12514 3049
rect 11480 3012 12204 3040
rect 11480 3000 11486 3012
rect 12176 2972 12204 3012
rect 12456 3009 12468 3043
rect 12502 3040 12514 3043
rect 12502 3012 12572 3040
rect 12502 3009 12514 3012
rect 12456 3003 12514 3009
rect 12544 2972 12572 3012
rect 12710 3000 12716 3052
rect 12768 3040 12774 3052
rect 13464 3049 13492 3080
rect 14829 3077 14841 3080
rect 14875 3077 14887 3111
rect 14829 3071 14887 3077
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 15804 3080 19104 3108
rect 15804 3068 15810 3080
rect 13449 3043 13507 3049
rect 12768 3012 12813 3040
rect 12912 3012 13308 3040
rect 12768 3000 12774 3012
rect 12912 2972 12940 3012
rect 9039 2944 12112 2972
rect 12176 2944 12940 2972
rect 13173 2975 13231 2981
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3694 2904 3700 2916
rect 2648 2876 3700 2904
rect 2648 2864 2654 2876
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 4249 2907 4307 2913
rect 4249 2873 4261 2907
rect 4295 2904 4307 2907
rect 5626 2904 5632 2916
rect 4295 2876 5632 2904
rect 4295 2873 4307 2876
rect 4249 2867 4307 2873
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 9861 2907 9919 2913
rect 9861 2873 9873 2907
rect 9907 2904 9919 2907
rect 11974 2904 11980 2916
rect 9907 2876 11980 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 1118 2796 1124 2848
rect 1176 2836 1182 2848
rect 1670 2836 1676 2848
rect 1176 2808 1676 2836
rect 1176 2796 1182 2808
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 2866 2836 2872 2848
rect 2827 2808 2872 2836
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 3568 2808 3617 2836
rect 3568 2796 3574 2808
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 3605 2799 3663 2805
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 6362 2836 6368 2848
rect 5583 2808 6368 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 9030 2836 9036 2848
rect 8435 2808 9036 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9398 2836 9404 2848
rect 9359 2808 9404 2836
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 11388 2808 11713 2836
rect 11388 2796 11394 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 12084 2836 12112 2944
rect 13173 2941 13185 2975
rect 13219 2941 13231 2975
rect 13280 2972 13308 3012
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3040 14703 3043
rect 14734 3040 14740 3052
rect 14691 3012 14740 3040
rect 14691 3009 14703 3012
rect 14645 3003 14703 3009
rect 14660 2972 14688 3003
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 14976 3012 15021 3040
rect 14976 3000 14982 3012
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15252 3012 16129 3040
rect 15252 3000 15258 3012
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 16117 3003 16175 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18966 3040 18972 3052
rect 17911 3012 18972 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 13280 2944 14688 2972
rect 13173 2935 13231 2941
rect 13188 2836 13216 2935
rect 17034 2932 17040 2984
rect 17092 2972 17098 2984
rect 17788 2972 17816 3003
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19076 3049 19104 3080
rect 19150 3068 19156 3120
rect 19208 3108 19214 3120
rect 26206 3108 26234 3148
rect 56965 3145 56977 3148
rect 57011 3145 57023 3179
rect 56965 3139 57023 3145
rect 19208 3080 26234 3108
rect 19208 3068 19214 3080
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 21266 3040 21272 3052
rect 21227 3012 21272 3040
rect 19705 3003 19763 3009
rect 17092 2944 17816 2972
rect 17092 2932 17098 2944
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 19720 2972 19748 3003
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23624 3012 23857 3040
rect 23624 3000 23630 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 23845 3003 23903 3009
rect 26206 3012 33701 3040
rect 18748 2944 19748 2972
rect 18748 2932 18754 2944
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 26206 2972 26234 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 33689 3003 33747 3009
rect 56686 3000 56692 3052
rect 56744 3040 56750 3052
rect 56781 3043 56839 3049
rect 56781 3040 56793 3043
rect 56744 3012 56793 3040
rect 56744 3000 56750 3012
rect 56781 3009 56793 3012
rect 56827 3009 56839 3043
rect 56781 3003 56839 3009
rect 20036 2944 26234 2972
rect 20036 2932 20042 2944
rect 33318 2932 33324 2984
rect 33376 2972 33382 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 33376 2944 33425 2972
rect 33376 2932 33382 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 17678 2904 17684 2916
rect 15979 2876 17684 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 17678 2864 17684 2876
rect 17736 2864 17742 2916
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 19521 2907 19579 2913
rect 19521 2904 19533 2907
rect 18012 2876 19533 2904
rect 18012 2864 18018 2876
rect 19521 2873 19533 2876
rect 19567 2873 19579 2907
rect 19521 2867 19579 2873
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 22186 2904 22192 2916
rect 21131 2876 22192 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 16666 2836 16672 2848
rect 12084 2808 16672 2836
rect 11701 2799 11759 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 16908 2808 16957 2836
rect 16908 2796 16914 2808
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 18877 2839 18935 2845
rect 18877 2805 18889 2839
rect 18923 2836 18935 2839
rect 19426 2836 19432 2848
rect 18923 2808 19432 2836
rect 18923 2805 18935 2808
rect 18877 2799 18935 2805
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 20441 2839 20499 2845
rect 20441 2836 20453 2839
rect 20220 2808 20453 2836
rect 20220 2796 20226 2808
rect 20441 2805 20453 2808
rect 20487 2805 20499 2839
rect 20441 2799 20499 2805
rect 21634 2796 21640 2848
rect 21692 2836 21698 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21692 2808 22017 2836
rect 21692 2796 21698 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 25096 2808 25329 2836
rect 25096 2796 25102 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 32585 2839 32643 2845
rect 32585 2836 32597 2839
rect 32364 2808 32597 2836
rect 32364 2796 32370 2808
rect 32585 2805 32597 2808
rect 32631 2805 32643 2839
rect 32585 2799 32643 2805
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35400 2808 35541 2836
rect 35400 2796 35406 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36780 2808 37473 2836
rect 36780 2796 36786 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 39945 2839 40003 2845
rect 39945 2836 39957 2839
rect 39724 2808 39957 2836
rect 39724 2796 39730 2808
rect 39945 2805 39957 2808
rect 39991 2805 40003 2839
rect 39945 2799 40003 2805
rect 42610 2796 42616 2848
rect 42668 2836 42674 2848
rect 42889 2839 42947 2845
rect 42889 2836 42901 2839
rect 42668 2808 42901 2836
rect 42668 2796 42674 2808
rect 42889 2805 42901 2808
rect 42935 2805 42947 2839
rect 42889 2799 42947 2805
rect 44082 2796 44088 2848
rect 44140 2836 44146 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 44140 2808 44373 2836
rect 44140 2796 44146 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 46934 2796 46940 2848
rect 46992 2836 46998 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 46992 2808 47777 2836
rect 46992 2796 46998 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 49878 2796 49884 2848
rect 49936 2836 49942 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49936 2808 50169 2836
rect 49936 2796 49942 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 52822 2796 52828 2848
rect 52880 2836 52886 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 52880 2808 53113 2836
rect 52880 2796 52886 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 54294 2796 54300 2848
rect 54352 2836 54358 2848
rect 54573 2839 54631 2845
rect 54573 2836 54585 2839
rect 54352 2808 54585 2836
rect 54352 2796 54358 2808
rect 54573 2805 54585 2808
rect 54619 2805 54631 2839
rect 54573 2799 54631 2805
rect 58161 2839 58219 2845
rect 58161 2805 58173 2839
rect 58207 2836 58219 2839
rect 58710 2836 58716 2848
rect 58207 2808 58716 2836
rect 58207 2805 58219 2808
rect 58161 2799 58219 2805
rect 58710 2796 58716 2808
rect 58768 2796 58774 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10284 2604 10425 2632
rect 10284 2592 10290 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14424 2604 18276 2632
rect 14424 2592 14430 2604
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 16117 2567 16175 2573
rect 5684 2536 10916 2564
rect 5684 2524 5690 2536
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6454 2496 6460 2508
rect 5859 2468 6460 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2428 3847 2431
rect 4706 2428 4712 2440
rect 3835 2400 4712 2428
rect 3835 2397 3847 2400
rect 3789 2391 3847 2397
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5534 2428 5540 2440
rect 5215 2400 5540 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6362 2428 6368 2440
rect 6323 2400 6368 2428
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8478 2428 8484 2440
rect 8435 2400 8484 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9030 2428 9036 2440
rect 8991 2400 9036 2428
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 10594 2428 10600 2440
rect 10555 2400 10600 2428
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10778 2428 10784 2440
rect 10739 2400 10784 2428
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10888 2437 10916 2536
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 17586 2564 17592 2576
rect 16163 2536 17592 2564
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 14461 2499 14519 2505
rect 14461 2465 14473 2499
rect 14507 2496 14519 2499
rect 15286 2496 15292 2508
rect 14507 2468 15292 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 16758 2496 16764 2508
rect 16719 2468 16764 2496
rect 16758 2456 16764 2468
rect 16816 2456 16822 2508
rect 17954 2496 17960 2508
rect 17236 2468 17960 2496
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2397 10931 2431
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 10873 2391 10931 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 14274 2428 14280 2440
rect 13587 2400 14280 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 14921 2391 14979 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17236 2437 17264 2468
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 18248 2496 18276 2604
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 25590 2632 25596 2644
rect 19116 2604 25452 2632
rect 25551 2604 25596 2632
rect 19116 2592 19122 2604
rect 18966 2524 18972 2576
rect 19024 2564 19030 2576
rect 21085 2567 21143 2573
rect 21085 2564 21097 2567
rect 19024 2536 21097 2564
rect 19024 2524 19030 2536
rect 21085 2533 21097 2536
rect 21131 2533 21143 2567
rect 21085 2527 21143 2533
rect 21174 2524 21180 2576
rect 21232 2564 21238 2576
rect 25314 2564 25320 2576
rect 21232 2536 25320 2564
rect 21232 2524 21238 2536
rect 25314 2524 25320 2536
rect 25372 2524 25378 2576
rect 25424 2564 25452 2604
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 25682 2592 25688 2644
rect 25740 2632 25746 2644
rect 27433 2635 27491 2641
rect 27433 2632 27445 2635
rect 25740 2604 27445 2632
rect 25740 2592 25746 2604
rect 27433 2601 27445 2604
rect 27479 2601 27491 2635
rect 28810 2632 28816 2644
rect 28771 2604 28816 2632
rect 27433 2595 27491 2601
rect 28810 2592 28816 2604
rect 28868 2592 28874 2644
rect 30282 2632 30288 2644
rect 30243 2604 30288 2632
rect 30282 2592 30288 2604
rect 30340 2592 30346 2644
rect 32355 2635 32413 2641
rect 32355 2632 32367 2635
rect 30392 2604 32367 2632
rect 30392 2564 30420 2604
rect 32355 2601 32367 2604
rect 32401 2601 32413 2635
rect 32355 2595 32413 2601
rect 37274 2592 37280 2644
rect 37332 2632 37338 2644
rect 45281 2635 45339 2641
rect 45281 2632 45293 2635
rect 37332 2604 45293 2632
rect 37332 2592 37338 2604
rect 45281 2601 45293 2604
rect 45327 2601 45339 2635
rect 45281 2595 45339 2601
rect 25424 2536 30420 2564
rect 30466 2524 30472 2576
rect 30524 2564 30530 2576
rect 54113 2567 54171 2573
rect 54113 2564 54125 2567
rect 30524 2536 54125 2564
rect 30524 2524 30530 2536
rect 54113 2533 54125 2536
rect 54159 2533 54171 2567
rect 54113 2527 54171 2533
rect 18248 2468 21404 2496
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17678 2428 17684 2440
rect 17639 2400 17684 2428
rect 17221 2391 17279 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 19150 2428 19156 2440
rect 18739 2400 19156 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19797 2431 19855 2437
rect 19797 2428 19809 2431
rect 19484 2400 19809 2428
rect 19484 2388 19490 2400
rect 19797 2397 19809 2400
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21140 2400 21281 2428
rect 21140 2388 21146 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21376 2428 21404 2468
rect 21450 2456 21456 2508
rect 21508 2496 21514 2508
rect 21508 2468 43024 2496
rect 21508 2456 21514 2468
rect 21542 2428 21548 2440
rect 21376 2400 21548 2428
rect 21269 2391 21327 2397
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 22186 2428 22192 2440
rect 22147 2400 22192 2428
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 23109 2431 23167 2437
rect 23109 2428 23121 2431
rect 22612 2400 23121 2428
rect 22612 2388 22618 2400
rect 23109 2397 23121 2400
rect 23155 2397 23167 2431
rect 23109 2391 23167 2397
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 24026 2428 24032 2440
rect 23891 2400 24032 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24670 2428 24676 2440
rect 24631 2400 24676 2428
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 25777 2431 25835 2437
rect 25777 2397 25789 2431
rect 25823 2428 25835 2431
rect 25958 2428 25964 2440
rect 25823 2400 25964 2428
rect 25823 2397 25835 2400
rect 25777 2391 25835 2397
rect 25958 2388 25964 2400
rect 26016 2388 26022 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 26510 2428 26516 2440
rect 26467 2400 26516 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 26510 2388 26516 2400
rect 26568 2388 26574 2440
rect 27430 2388 27436 2440
rect 27488 2428 27494 2440
rect 27617 2431 27675 2437
rect 27617 2428 27629 2431
rect 27488 2400 27629 2428
rect 27488 2388 27494 2400
rect 27617 2397 27629 2400
rect 27663 2397 27675 2431
rect 27617 2391 27675 2397
rect 27982 2388 27988 2440
rect 28040 2428 28046 2440
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 28040 2400 28273 2428
rect 28040 2388 28046 2400
rect 28261 2397 28273 2400
rect 28307 2397 28319 2431
rect 28261 2391 28319 2397
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 28960 2400 29009 2428
rect 28960 2388 28966 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 28997 2391 29055 2397
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29512 2400 29745 2428
rect 29512 2388 29518 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30374 2388 30380 2440
rect 30432 2428 30438 2440
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 30432 2400 30481 2428
rect 30432 2388 30438 2400
rect 30469 2397 30481 2400
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 30892 2400 31125 2428
rect 30892 2388 30898 2400
rect 31113 2397 31125 2400
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 31846 2388 31852 2440
rect 31904 2428 31910 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31904 2400 32137 2428
rect 31904 2388 31910 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34057 2431 34115 2437
rect 34057 2428 34069 2431
rect 33836 2400 34069 2428
rect 33836 2388 33842 2400
rect 34057 2397 34069 2400
rect 34103 2397 34115 2431
rect 34057 2391 34115 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 35158 2428 35164 2440
rect 35119 2400 35164 2428
rect 34885 2391 34943 2397
rect 35158 2388 35164 2400
rect 35216 2388 35222 2440
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 35866 2400 38117 2428
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 9815 2332 10916 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10888 2304 10916 2332
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 21174 2360 21180 2372
rect 15988 2332 21180 2360
rect 15988 2320 15994 2332
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 35866 2360 35894 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38194 2388 38200 2440
rect 38252 2428 38258 2440
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38252 2400 38761 2428
rect 38252 2388 38258 2400
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 39132 2400 41184 2428
rect 21468 2332 35894 2360
rect 3050 2252 3056 2304
rect 3108 2292 3114 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3108 2264 3985 2292
rect 3108 2252 3114 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6549 2295 6607 2301
rect 6549 2292 6561 2295
rect 6052 2264 6561 2292
rect 6052 2252 6058 2264
rect 6549 2261 6561 2264
rect 6595 2261 6607 2295
rect 6549 2255 6607 2261
rect 7561 2295 7619 2301
rect 7561 2261 7573 2295
rect 7607 2292 7619 2295
rect 7926 2292 7932 2304
rect 7607 2264 7932 2292
rect 7607 2261 7619 2264
rect 7561 2255 7619 2261
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 8996 2264 9229 2292
rect 8996 2252 9002 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 10870 2252 10876 2304
rect 10928 2252 10934 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 11940 2264 12173 2292
rect 11940 2252 11946 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12161 2255 12219 2261
rect 12713 2295 12771 2301
rect 12713 2261 12725 2295
rect 12759 2292 12771 2295
rect 13814 2292 13820 2304
rect 12759 2264 13820 2292
rect 12759 2261 12771 2264
rect 12713 2255 12771 2261
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15105 2295 15163 2301
rect 15105 2292 15117 2295
rect 14884 2264 15117 2292
rect 14884 2252 14890 2264
rect 15105 2261 15117 2264
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17276 2264 17877 2292
rect 17276 2252 17282 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 19978 2292 19984 2304
rect 19939 2264 19984 2292
rect 17865 2255 17923 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 21468 2292 21496 2332
rect 36262 2320 36268 2372
rect 36320 2360 36326 2372
rect 36449 2363 36507 2369
rect 36449 2360 36461 2363
rect 36320 2332 36461 2360
rect 36320 2320 36326 2332
rect 36449 2329 36461 2332
rect 36495 2329 36507 2363
rect 36449 2323 36507 2329
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 37921 2363 37979 2369
rect 37921 2360 37933 2363
rect 37792 2332 37933 2360
rect 37792 2320 37798 2332
rect 37921 2329 37933 2332
rect 37967 2329 37979 2363
rect 37921 2323 37979 2329
rect 38562 2320 38568 2372
rect 38620 2360 38626 2372
rect 39132 2360 39160 2400
rect 38620 2332 39160 2360
rect 38620 2320 38626 2332
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 39264 2332 40325 2360
rect 39264 2320 39270 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 41032 2363 41090 2369
rect 41032 2360 41044 2363
rect 40644 2332 41044 2360
rect 40644 2320 40650 2332
rect 41032 2329 41044 2332
rect 41078 2329 41090 2363
rect 41156 2360 41184 2400
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 41877 2431 41935 2437
rect 41877 2428 41889 2431
rect 41380 2400 41889 2428
rect 41380 2388 41386 2400
rect 41877 2397 41889 2400
rect 41923 2397 41935 2431
rect 41877 2391 41935 2397
rect 41156 2332 41276 2360
rect 41032 2323 41090 2329
rect 20128 2264 21496 2292
rect 20128 2252 20134 2264
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 22373 2295 22431 2301
rect 22373 2292 22385 2295
rect 22152 2264 22385 2292
rect 22152 2252 22158 2264
rect 22373 2261 22385 2264
rect 22419 2261 22431 2295
rect 22373 2255 22431 2261
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 24857 2295 24915 2301
rect 24857 2292 24869 2295
rect 24636 2264 24869 2292
rect 24636 2252 24642 2264
rect 24857 2261 24869 2264
rect 24903 2261 24915 2295
rect 24857 2255 24915 2261
rect 25314 2252 25320 2304
rect 25372 2292 25378 2304
rect 36541 2295 36599 2301
rect 36541 2292 36553 2295
rect 25372 2264 36553 2292
rect 25372 2252 25378 2264
rect 36541 2261 36553 2264
rect 36587 2261 36599 2295
rect 40402 2292 40408 2304
rect 40363 2264 40408 2292
rect 36541 2255 36599 2261
rect 40402 2252 40408 2264
rect 40460 2252 40466 2304
rect 40494 2252 40500 2304
rect 40552 2292 40558 2304
rect 41141 2295 41199 2301
rect 41141 2292 41153 2295
rect 40552 2264 41153 2292
rect 40552 2252 40558 2264
rect 41141 2261 41153 2264
rect 41187 2261 41199 2295
rect 41248 2292 41276 2332
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 42116 2332 42901 2360
rect 42116 2320 42122 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42996 2360 43024 2468
rect 43070 2388 43076 2440
rect 43128 2428 43134 2440
rect 43128 2400 43173 2428
rect 43128 2388 43134 2400
rect 43530 2388 43536 2440
rect 43588 2428 43594 2440
rect 43625 2431 43683 2437
rect 43625 2428 43637 2431
rect 43588 2400 43637 2428
rect 43588 2388 43594 2400
rect 43625 2397 43637 2400
rect 43671 2397 43683 2431
rect 43625 2391 43683 2397
rect 45002 2388 45008 2440
rect 45060 2428 45066 2440
rect 45097 2431 45155 2437
rect 45097 2428 45109 2431
rect 45060 2400 45109 2428
rect 45060 2388 45066 2400
rect 45097 2397 45109 2400
rect 45143 2397 45155 2431
rect 45097 2391 45155 2397
rect 45462 2388 45468 2440
rect 45520 2428 45526 2440
rect 46017 2431 46075 2437
rect 46017 2428 46029 2431
rect 45520 2400 46029 2428
rect 45520 2388 45526 2400
rect 46017 2397 46029 2400
rect 46063 2397 46075 2431
rect 46017 2391 46075 2397
rect 46474 2388 46480 2440
rect 46532 2428 46538 2440
rect 46569 2431 46627 2437
rect 46569 2428 46581 2431
rect 46532 2400 46581 2428
rect 46532 2388 46538 2400
rect 46569 2397 46581 2400
rect 46615 2397 46627 2431
rect 46569 2391 46627 2397
rect 47946 2388 47952 2440
rect 48004 2428 48010 2440
rect 48041 2431 48099 2437
rect 48041 2428 48053 2431
rect 48004 2400 48053 2428
rect 48004 2388 48010 2400
rect 48041 2397 48053 2400
rect 48087 2397 48099 2431
rect 48041 2391 48099 2397
rect 48406 2388 48412 2440
rect 48464 2428 48470 2440
rect 48961 2431 49019 2437
rect 48961 2428 48973 2431
rect 48464 2400 48973 2428
rect 48464 2388 48470 2400
rect 48961 2397 48973 2400
rect 49007 2397 49019 2431
rect 48961 2391 49019 2397
rect 49418 2388 49424 2440
rect 49476 2428 49482 2440
rect 50157 2431 50215 2437
rect 50157 2428 50169 2431
rect 49476 2400 50169 2428
rect 49476 2388 49482 2400
rect 50157 2397 50169 2400
rect 50203 2397 50215 2431
rect 50157 2391 50215 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 50985 2431 51043 2437
rect 50985 2428 50997 2431
rect 50948 2400 50997 2428
rect 50948 2388 50954 2400
rect 50985 2397 50997 2400
rect 51031 2397 51043 2431
rect 50985 2391 51043 2397
rect 51350 2388 51356 2440
rect 51408 2428 51414 2440
rect 51905 2431 51963 2437
rect 51905 2428 51917 2431
rect 51408 2400 51917 2428
rect 51408 2388 51414 2400
rect 51905 2397 51917 2400
rect 51951 2397 51963 2431
rect 51905 2391 51963 2397
rect 52362 2388 52368 2440
rect 52420 2428 52426 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52420 2400 52745 2428
rect 52420 2388 52426 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53834 2388 53840 2440
rect 53892 2428 53898 2440
rect 53929 2431 53987 2437
rect 53929 2428 53941 2431
rect 53892 2400 53941 2428
rect 53892 2388 53898 2400
rect 53929 2397 53941 2400
rect 53975 2397 53987 2431
rect 53929 2391 53987 2397
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 55272 2400 55321 2428
rect 55272 2388 55278 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 55766 2388 55772 2440
rect 55824 2428 55830 2440
rect 56229 2431 56287 2437
rect 56229 2428 56241 2431
rect 55824 2400 56241 2428
rect 55824 2388 55830 2400
rect 56229 2397 56241 2400
rect 56275 2397 56287 2431
rect 56229 2391 56287 2397
rect 57238 2388 57244 2440
rect 57296 2428 57302 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 57296 2400 58081 2428
rect 57296 2388 57302 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 56965 2363 57023 2369
rect 42996 2332 48268 2360
rect 42889 2323 42947 2329
rect 43809 2295 43867 2301
rect 43809 2292 43821 2295
rect 41248 2264 43821 2292
rect 41141 2255 41199 2261
rect 43809 2261 43821 2264
rect 43855 2261 43867 2295
rect 46750 2292 46756 2304
rect 46711 2264 46756 2292
rect 43809 2255 43867 2261
rect 46750 2252 46756 2264
rect 46808 2252 46814 2304
rect 48240 2301 48268 2332
rect 56965 2329 56977 2363
rect 57011 2360 57023 2363
rect 58158 2360 58164 2372
rect 57011 2332 58164 2360
rect 57011 2329 57023 2332
rect 56965 2323 57023 2329
rect 58158 2320 58164 2332
rect 58216 2320 58222 2372
rect 48225 2295 48283 2301
rect 48225 2261 48237 2295
rect 48271 2261 48283 2295
rect 48225 2255 48283 2261
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 50341 2295 50399 2301
rect 50341 2292 50353 2295
rect 48372 2264 50353 2292
rect 48372 2252 48378 2264
rect 50341 2261 50353 2264
rect 50387 2261 50399 2295
rect 51166 2292 51172 2304
rect 51127 2264 51172 2292
rect 50341 2255 50399 2261
rect 51166 2252 51172 2264
rect 51224 2252 51230 2304
rect 52914 2292 52920 2304
rect 52875 2264 52920 2292
rect 52914 2252 52920 2264
rect 52972 2252 52978 2304
rect 55490 2292 55496 2304
rect 55451 2264 55496 2292
rect 55490 2252 55496 2264
rect 55548 2252 55554 2304
rect 57054 2292 57060 2304
rect 57015 2264 57060 2292
rect 57054 2252 57060 2264
rect 57112 2252 57118 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 21450 2088 21456 2100
rect 14608 2060 21456 2088
rect 14608 2048 14614 2060
rect 21450 2048 21456 2060
rect 21508 2048 21514 2100
rect 21542 2048 21548 2100
rect 21600 2088 21606 2100
rect 46750 2088 46756 2100
rect 21600 2060 46756 2088
rect 21600 2048 21606 2060
rect 46750 2048 46756 2060
rect 46808 2048 46814 2100
rect 15654 1980 15660 2032
rect 15712 2020 15718 2032
rect 20070 2020 20076 2032
rect 15712 1992 20076 2020
rect 15712 1980 15718 1992
rect 20070 1980 20076 1992
rect 20128 1980 20134 2032
rect 20806 1980 20812 2032
rect 20864 2020 20870 2032
rect 51166 2020 51172 2032
rect 20864 1992 51172 2020
rect 20864 1980 20870 1992
rect 51166 1980 51172 1992
rect 51224 1980 51230 2032
rect 15010 1912 15016 1964
rect 15068 1952 15074 1964
rect 43070 1952 43076 1964
rect 15068 1924 43076 1952
rect 15068 1912 15074 1924
rect 43070 1912 43076 1924
rect 43128 1912 43134 1964
rect 15102 1844 15108 1896
rect 15160 1884 15166 1896
rect 40402 1884 40408 1896
rect 15160 1856 40408 1884
rect 15160 1844 15166 1856
rect 40402 1844 40408 1856
rect 40460 1844 40466 1896
rect 20622 1776 20628 1828
rect 20680 1816 20686 1828
rect 30466 1816 30472 1828
rect 20680 1788 30472 1816
rect 20680 1776 20686 1788
rect 30466 1776 30472 1788
rect 30524 1776 30530 1828
rect 17310 1708 17316 1760
rect 17368 1748 17374 1760
rect 57054 1748 57060 1760
rect 17368 1720 57060 1748
rect 17368 1708 17374 1720
rect 57054 1708 57060 1720
rect 57112 1708 57118 1760
rect 20530 1640 20536 1692
rect 20588 1680 20594 1692
rect 55490 1680 55496 1692
rect 20588 1652 55496 1680
rect 20588 1640 20594 1652
rect 55490 1640 55496 1652
rect 55548 1640 55554 1692
rect 15838 1572 15844 1624
rect 15896 1612 15902 1624
rect 35158 1612 35164 1624
rect 15896 1584 35164 1612
rect 15896 1572 15902 1584
rect 35158 1572 35164 1584
rect 35216 1572 35222 1624
rect 20438 1504 20444 1556
rect 20496 1544 20502 1556
rect 52914 1544 52920 1556
rect 20496 1516 52920 1544
rect 20496 1504 20502 1516
rect 52914 1504 52920 1516
rect 52972 1504 52978 1556
rect 2774 1436 2780 1488
rect 2832 1476 2838 1488
rect 5166 1476 5172 1488
rect 2832 1448 5172 1476
rect 2832 1436 2838 1448
rect 5166 1436 5172 1448
rect 5224 1436 5230 1488
rect 19242 1436 19248 1488
rect 19300 1476 19306 1488
rect 48314 1476 48320 1488
rect 19300 1448 48320 1476
rect 19300 1436 19306 1448
rect 48314 1436 48320 1448
rect 48372 1436 48378 1488
rect 16022 1368 16028 1420
rect 16080 1408 16086 1420
rect 40494 1408 40500 1420
rect 16080 1380 40500 1408
rect 16080 1368 16086 1380
rect 40494 1368 40500 1380
rect 40552 1368 40558 1420
rect 3418 1164 3424 1216
rect 3476 1204 3482 1216
rect 7098 1204 7104 1216
rect 3476 1176 7104 1204
rect 3476 1164 3482 1176
rect 7098 1164 7104 1176
rect 7156 1164 7162 1216
<< via1 >>
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1584 39627 1636 39636
rect 1584 39593 1593 39627
rect 1593 39593 1627 39627
rect 1627 39593 1636 39627
rect 1584 39584 1636 39593
rect 2780 39584 2832 39636
rect 3700 39584 3752 39636
rect 26240 39584 26292 39636
rect 41420 39627 41472 39636
rect 41420 39593 41429 39627
rect 41429 39593 41463 39627
rect 41463 39593 41472 39627
rect 41420 39584 41472 39593
rect 48688 39584 48740 39636
rect 56140 39584 56192 39636
rect 18696 39448 18748 39500
rect 2136 39423 2188 39432
rect 2136 39389 2145 39423
rect 2145 39389 2179 39423
rect 2179 39389 2188 39423
rect 2136 39380 2188 39389
rect 6644 39380 6696 39432
rect 2320 39312 2372 39364
rect 3056 39287 3108 39296
rect 3056 39253 3065 39287
rect 3065 39253 3099 39287
rect 3099 39253 3108 39287
rect 3056 39244 3108 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 2504 38904 2556 38956
rect 1584 38743 1636 38752
rect 1584 38709 1593 38743
rect 1593 38709 1627 38743
rect 1627 38709 1636 38743
rect 1584 38700 1636 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1492 38496 1544 38548
rect 1492 38292 1544 38344
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 1676 37816 1728 37868
rect 1584 37655 1636 37664
rect 1584 37621 1593 37655
rect 1593 37621 1627 37655
rect 1627 37621 1636 37655
rect 1584 37612 1636 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 1768 36728 1820 36780
rect 1584 36635 1636 36644
rect 1584 36601 1593 36635
rect 1593 36601 1627 36635
rect 1627 36601 1636 36635
rect 1584 36592 1636 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1860 36116 1912 36168
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1952 35028 2004 35080
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 2872 34688 2924 34740
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6276 33940 6328 33992
rect 1584 33847 1636 33856
rect 1584 33813 1593 33847
rect 1593 33813 1627 33847
rect 1627 33813 1636 33847
rect 1584 33804 1636 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 1584 33507 1636 33516
rect 1584 33473 1593 33507
rect 1593 33473 1627 33507
rect 1627 33473 1636 33507
rect 1584 33464 1636 33473
rect 2412 33507 2464 33516
rect 2412 33473 2421 33507
rect 2421 33473 2455 33507
rect 2455 33473 2464 33507
rect 2412 33464 2464 33473
rect 4988 33328 5040 33380
rect 2136 33260 2188 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4620 32988 4672 33040
rect 4988 32963 5040 32972
rect 4988 32929 4997 32963
rect 4997 32929 5031 32963
rect 5031 32929 5040 32963
rect 4988 32920 5040 32929
rect 5080 32963 5132 32972
rect 5080 32929 5089 32963
rect 5089 32929 5123 32963
rect 5123 32929 5132 32963
rect 5080 32920 5132 32929
rect 2136 32895 2188 32904
rect 2136 32861 2170 32895
rect 2170 32861 2188 32895
rect 2136 32852 2188 32861
rect 2780 32784 2832 32836
rect 4804 32716 4856 32768
rect 4896 32759 4948 32768
rect 4896 32725 4905 32759
rect 4905 32725 4939 32759
rect 4939 32725 4948 32759
rect 4896 32716 4948 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 1584 32555 1636 32564
rect 1584 32521 1593 32555
rect 1593 32521 1627 32555
rect 1627 32521 1636 32555
rect 1584 32512 1636 32521
rect 2412 32555 2464 32564
rect 2412 32521 2421 32555
rect 2421 32521 2455 32555
rect 2455 32521 2464 32555
rect 2412 32512 2464 32521
rect 2872 32555 2924 32564
rect 2872 32521 2881 32555
rect 2881 32521 2915 32555
rect 2915 32521 2924 32555
rect 2872 32512 2924 32521
rect 4896 32512 4948 32564
rect 4620 32444 4672 32496
rect 4712 32419 4764 32428
rect 4712 32385 4746 32419
rect 4746 32385 4764 32419
rect 4712 32376 4764 32385
rect 3148 32308 3200 32360
rect 2780 32240 2832 32292
rect 7564 32172 7616 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4712 31968 4764 32020
rect 2964 31900 3016 31952
rect 1584 31807 1636 31816
rect 1584 31773 1593 31807
rect 1593 31773 1627 31807
rect 1627 31773 1636 31807
rect 1584 31764 1636 31773
rect 3056 31807 3108 31816
rect 3056 31773 3065 31807
rect 3065 31773 3099 31807
rect 3099 31773 3108 31807
rect 3056 31764 3108 31773
rect 4804 31764 4856 31816
rect 2872 31671 2924 31680
rect 2872 31637 2881 31671
rect 2881 31637 2915 31671
rect 2915 31637 2924 31671
rect 2872 31628 2924 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2872 31356 2924 31408
rect 4620 31356 4672 31408
rect 3424 31288 3476 31340
rect 4896 31331 4948 31340
rect 4896 31297 4905 31331
rect 4905 31297 4939 31331
rect 4939 31297 4948 31331
rect 4896 31288 4948 31297
rect 4988 31331 5040 31340
rect 4988 31297 4997 31331
rect 4997 31297 5031 31331
rect 5031 31297 5040 31331
rect 4988 31288 5040 31297
rect 2780 31220 2832 31272
rect 1584 31195 1636 31204
rect 1584 31161 1593 31195
rect 1593 31161 1627 31195
rect 1627 31161 1636 31195
rect 1584 31152 1636 31161
rect 4620 31152 4672 31204
rect 2872 31084 2924 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3056 30880 3108 30932
rect 2964 30787 3016 30796
rect 2964 30753 2973 30787
rect 2973 30753 3007 30787
rect 3007 30753 3016 30787
rect 2964 30744 3016 30753
rect 3148 30787 3200 30796
rect 3148 30753 3157 30787
rect 3157 30753 3191 30787
rect 3191 30753 3200 30787
rect 3148 30744 3200 30753
rect 4896 30744 4948 30796
rect 5080 30744 5132 30796
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 2872 30719 2924 30728
rect 2872 30685 2881 30719
rect 2881 30685 2915 30719
rect 2915 30685 2924 30719
rect 2872 30676 2924 30685
rect 4712 30540 4764 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4988 30336 5040 30388
rect 7748 30268 7800 30320
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 2780 30064 2832 30116
rect 2964 30064 3016 30116
rect 1584 30039 1636 30048
rect 1584 30005 1593 30039
rect 1593 30005 1627 30039
rect 1627 30005 1636 30039
rect 1584 29996 1636 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2688 29792 2740 29844
rect 4896 29656 4948 29708
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 4988 29588 5040 29640
rect 4712 29520 4764 29572
rect 2872 29452 2924 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2872 29291 2924 29300
rect 2872 29257 2881 29291
rect 2881 29257 2915 29291
rect 2915 29257 2924 29291
rect 2872 29248 2924 29257
rect 7656 29180 7708 29232
rect 2780 29155 2832 29164
rect 2780 29121 2789 29155
rect 2789 29121 2823 29155
rect 2823 29121 2832 29155
rect 2780 29112 2832 29121
rect 2688 29044 2740 29096
rect 1584 29019 1636 29028
rect 1584 28985 1593 29019
rect 1593 28985 1627 29019
rect 1627 28985 1636 29019
rect 1584 28976 1636 28985
rect 2504 28908 2556 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2964 28500 3016 28552
rect 2320 28432 2372 28484
rect 2780 28364 2832 28416
rect 3792 28364 3844 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2320 28203 2372 28212
rect 2320 28169 2329 28203
rect 2329 28169 2363 28203
rect 2363 28169 2372 28203
rect 2320 28160 2372 28169
rect 1400 28024 1452 28076
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 2596 28024 2648 28076
rect 3884 28067 3936 28076
rect 3884 28033 3893 28067
rect 3893 28033 3927 28067
rect 3927 28033 3936 28067
rect 3884 28024 3936 28033
rect 2504 27888 2556 27940
rect 2688 27956 2740 28008
rect 3976 27999 4028 28008
rect 3976 27965 3985 27999
rect 3985 27965 4019 27999
rect 4019 27965 4028 27999
rect 3976 27956 4028 27965
rect 2688 27820 2740 27872
rect 4068 27820 4120 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3976 27616 4028 27668
rect 2320 27412 2372 27464
rect 3056 27455 3108 27464
rect 3056 27421 3065 27455
rect 3065 27421 3099 27455
rect 3099 27421 3108 27455
rect 3056 27412 3108 27421
rect 2964 27344 3016 27396
rect 3700 27412 3752 27464
rect 13084 27412 13136 27464
rect 3976 27344 4028 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 2228 27319 2280 27328
rect 2228 27285 2237 27319
rect 2237 27285 2271 27319
rect 2271 27285 2280 27319
rect 2228 27276 2280 27285
rect 3884 27276 3936 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 3976 27115 4028 27124
rect 3976 27081 3985 27115
rect 3985 27081 4019 27115
rect 4019 27081 4028 27115
rect 3976 27072 4028 27081
rect 2228 27004 2280 27056
rect 2964 26936 3016 26988
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 3148 26775 3200 26784
rect 3148 26741 3157 26775
rect 3157 26741 3191 26775
rect 3191 26741 3200 26775
rect 3148 26732 3200 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2320 26528 2372 26580
rect 3148 26528 3200 26580
rect 2688 26435 2740 26444
rect 2688 26401 2697 26435
rect 2697 26401 2731 26435
rect 2731 26401 2740 26435
rect 2688 26392 2740 26401
rect 2872 26435 2924 26444
rect 2872 26401 2881 26435
rect 2881 26401 2915 26435
rect 2915 26401 2924 26435
rect 3884 26435 3936 26444
rect 2872 26392 2924 26401
rect 3884 26401 3893 26435
rect 3893 26401 3927 26435
rect 3927 26401 3936 26435
rect 3884 26392 3936 26401
rect 4712 26460 4764 26512
rect 15752 26392 15804 26444
rect 3976 26324 4028 26376
rect 3148 26256 3200 26308
rect 3792 26299 3844 26308
rect 3792 26265 3801 26299
rect 3801 26265 3835 26299
rect 3835 26265 3844 26299
rect 3792 26256 3844 26265
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 3884 25891 3936 25900
rect 3884 25857 3893 25891
rect 3893 25857 3927 25891
rect 3927 25857 3936 25891
rect 3884 25848 3936 25857
rect 3608 25644 3660 25696
rect 4068 25644 4120 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3976 25440 4028 25492
rect 2780 25236 2832 25288
rect 3700 25236 3752 25288
rect 12256 25236 12308 25288
rect 4068 25211 4120 25220
rect 4068 25177 4102 25211
rect 4102 25177 4120 25211
rect 4068 25168 4120 25177
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3884 24896 3936 24948
rect 3976 24828 4028 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 2228 24760 2280 24812
rect 3608 24760 3660 24812
rect 2596 24692 2648 24744
rect 2688 24624 2740 24676
rect 2136 24556 2188 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2136 24191 2188 24200
rect 2136 24157 2170 24191
rect 2170 24157 2188 24191
rect 2136 24148 2188 24157
rect 2780 24080 2832 24132
rect 1400 24012 1452 24064
rect 1768 24012 1820 24064
rect 1860 24012 1912 24064
rect 2136 24012 2188 24064
rect 3332 24012 3384 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 2228 23851 2280 23860
rect 2228 23817 2237 23851
rect 2237 23817 2271 23851
rect 2271 23817 2280 23851
rect 2228 23808 2280 23817
rect 2688 23851 2740 23860
rect 2688 23817 2697 23851
rect 2697 23817 2731 23851
rect 2731 23817 2740 23851
rect 2688 23808 2740 23817
rect 1860 23672 1912 23724
rect 3332 23672 3384 23724
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 2688 23604 2740 23656
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 2780 23060 2832 23112
rect 4068 23060 4120 23112
rect 4620 22992 4672 23044
rect 3884 22924 3936 22976
rect 3976 22924 4028 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1492 22720 1544 22772
rect 1952 22720 2004 22772
rect 3884 22763 3936 22772
rect 3884 22729 3893 22763
rect 3893 22729 3927 22763
rect 3927 22729 3936 22763
rect 3884 22720 3936 22729
rect 4620 22763 4672 22772
rect 4620 22729 4629 22763
rect 4629 22729 4663 22763
rect 4663 22729 4672 22763
rect 4620 22720 4672 22729
rect 3700 22652 3752 22704
rect 3976 22652 4028 22704
rect 1492 22584 1544 22636
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 2596 22516 2648 22568
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 2136 22380 2188 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5448 22176 5500 22228
rect 4068 22108 4120 22160
rect 4712 22040 4764 22092
rect 2136 22015 2188 22024
rect 2136 21981 2170 22015
rect 2170 21981 2188 22015
rect 2136 21972 2188 21981
rect 3976 21972 4028 22024
rect 6184 21972 6236 22024
rect 9680 21972 9732 22024
rect 2780 21904 2832 21956
rect 4804 21904 4856 21956
rect 8024 21904 8076 21956
rect 3240 21879 3292 21888
rect 3240 21845 3249 21879
rect 3249 21845 3283 21879
rect 3283 21845 3292 21879
rect 3240 21836 3292 21845
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 6276 21836 6328 21888
rect 8116 21836 8168 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2412 21632 2464 21684
rect 3976 21675 4028 21684
rect 3976 21641 3985 21675
rect 3985 21641 4019 21675
rect 4019 21641 4028 21675
rect 3976 21632 4028 21641
rect 17316 21564 17368 21616
rect 2688 21471 2740 21480
rect 2688 21437 2697 21471
rect 2697 21437 2731 21471
rect 2731 21437 2740 21471
rect 2688 21428 2740 21437
rect 2596 21360 2648 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 3240 21496 3292 21548
rect 3332 21496 3384 21548
rect 3700 21539 3752 21548
rect 3700 21505 3709 21539
rect 3709 21505 3743 21539
rect 3743 21505 3752 21539
rect 3700 21496 3752 21505
rect 3792 21539 3844 21548
rect 3792 21505 3801 21539
rect 3801 21505 3835 21539
rect 3835 21505 3844 21539
rect 3792 21496 3844 21505
rect 9680 21496 9732 21548
rect 10416 21496 10468 21548
rect 10968 21335 11020 21344
rect 10968 21301 10977 21335
rect 10977 21301 11011 21335
rect 11011 21301 11020 21335
rect 10968 21292 11020 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2688 21088 2740 21140
rect 7564 21131 7616 21140
rect 7564 21097 7573 21131
rect 7573 21097 7607 21131
rect 7607 21097 7616 21131
rect 7564 21088 7616 21097
rect 9404 21131 9456 21140
rect 9404 21097 9413 21131
rect 9413 21097 9447 21131
rect 9447 21097 9456 21131
rect 9404 21088 9456 21097
rect 10416 21131 10468 21140
rect 10416 21097 10425 21131
rect 10425 21097 10459 21131
rect 10459 21097 10468 21131
rect 10416 21088 10468 21097
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 7748 21020 7800 21072
rect 4712 20952 4764 21004
rect 6184 20995 6236 21004
rect 6184 20961 6193 20995
rect 6193 20961 6227 20995
rect 6227 20961 6236 20995
rect 6184 20952 6236 20961
rect 8116 20995 8168 21004
rect 8116 20961 8125 20995
rect 8125 20961 8159 20995
rect 8159 20961 8168 20995
rect 8116 20952 8168 20961
rect 10968 21020 11020 21072
rect 9956 20952 10008 21004
rect 1400 20884 1452 20936
rect 2412 20927 2464 20936
rect 2412 20893 2421 20927
rect 2421 20893 2455 20927
rect 2455 20893 2464 20927
rect 2412 20884 2464 20893
rect 8300 20884 8352 20936
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10968 20884 11020 20936
rect 4712 20816 4764 20868
rect 7104 20816 7156 20868
rect 12532 20884 12584 20936
rect 12440 20816 12492 20868
rect 2228 20791 2280 20800
rect 2228 20757 2237 20791
rect 2237 20757 2271 20791
rect 2271 20757 2280 20791
rect 2228 20748 2280 20757
rect 8392 20791 8444 20800
rect 8392 20757 8401 20791
rect 8401 20757 8435 20791
rect 8435 20757 8444 20791
rect 8392 20748 8444 20757
rect 10968 20748 11020 20800
rect 14648 20859 14700 20868
rect 14648 20825 14682 20859
rect 14682 20825 14700 20859
rect 14648 20816 14700 20825
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 3792 20544 3844 20596
rect 7104 20587 7156 20596
rect 7104 20553 7113 20587
rect 7113 20553 7147 20587
rect 7147 20553 7156 20587
rect 7104 20544 7156 20553
rect 7472 20544 7524 20596
rect 8024 20587 8076 20596
rect 2228 20519 2280 20528
rect 2228 20485 2262 20519
rect 2262 20485 2280 20519
rect 2228 20476 2280 20485
rect 2780 20408 2832 20460
rect 8024 20553 8033 20587
rect 8033 20553 8067 20587
rect 8067 20553 8076 20587
rect 8024 20544 8076 20553
rect 8392 20587 8444 20596
rect 8392 20553 8401 20587
rect 8401 20553 8435 20587
rect 8435 20553 8444 20587
rect 8392 20544 8444 20553
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 14648 20587 14700 20596
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 7840 20340 7892 20392
rect 7656 20272 7708 20324
rect 8576 20408 8628 20460
rect 12532 20408 12584 20460
rect 12716 20408 12768 20460
rect 13544 20408 13596 20460
rect 15016 20451 15068 20460
rect 15016 20417 15025 20451
rect 15025 20417 15059 20451
rect 15059 20417 15068 20451
rect 15016 20408 15068 20417
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2412 20000 2464 20052
rect 7840 20043 7892 20052
rect 1584 19975 1636 19984
rect 1584 19941 1593 19975
rect 1593 19941 1627 19975
rect 1627 19941 1636 19975
rect 1584 19932 1636 19941
rect 7840 20009 7849 20043
rect 7849 20009 7883 20043
rect 7883 20009 7892 20043
rect 7840 20000 7892 20009
rect 12716 20043 12768 20052
rect 9404 19932 9456 19984
rect 12716 20009 12725 20043
rect 12725 20009 12759 20043
rect 12759 20009 12768 20043
rect 12716 20000 12768 20009
rect 15016 20043 15068 20052
rect 12808 19932 12860 19984
rect 15016 20009 15025 20043
rect 15025 20009 15059 20043
rect 15059 20009 15068 20043
rect 15016 20000 15068 20009
rect 2136 19864 2188 19916
rect 2412 19864 2464 19916
rect 2596 19864 2648 19916
rect 7564 19907 7616 19916
rect 7564 19873 7573 19907
rect 7573 19873 7607 19907
rect 7607 19873 7616 19907
rect 7564 19864 7616 19873
rect 3332 19728 3384 19780
rect 8300 19796 8352 19848
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 13084 19796 13136 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15752 19796 15804 19848
rect 18052 19728 18104 19780
rect 2688 19703 2740 19712
rect 2688 19669 2697 19703
rect 2697 19669 2731 19703
rect 2731 19669 2740 19703
rect 2688 19660 2740 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2688 19456 2740 19508
rect 3424 19456 3476 19508
rect 1400 19320 1452 19372
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 2780 19320 2832 19372
rect 4068 19320 4120 19372
rect 7104 19388 7156 19440
rect 7656 19320 7708 19372
rect 12532 19388 12584 19440
rect 8300 19363 8352 19372
rect 8300 19329 8309 19363
rect 8309 19329 8343 19363
rect 8343 19329 8352 19363
rect 8300 19320 8352 19329
rect 9404 19363 9456 19372
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 12348 19320 12400 19372
rect 14280 19320 14332 19372
rect 14648 19320 14700 19372
rect 15200 19388 15252 19440
rect 2688 19116 2740 19168
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 9680 19252 9732 19304
rect 12900 19295 12952 19304
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 12900 19252 12952 19261
rect 12256 19184 12308 19236
rect 16856 19252 16908 19304
rect 9772 19116 9824 19168
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 13176 19159 13228 19168
rect 13176 19125 13185 19159
rect 13185 19125 13219 19159
rect 13219 19125 13228 19159
rect 13176 19116 13228 19125
rect 13728 19116 13780 19168
rect 15568 19116 15620 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1860 18912 1912 18964
rect 1768 18776 1820 18828
rect 2228 18708 2280 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 8392 18844 8444 18896
rect 7748 18776 7800 18828
rect 12808 18912 12860 18964
rect 13728 18912 13780 18964
rect 16856 18955 16908 18964
rect 16856 18921 16865 18955
rect 16865 18921 16899 18955
rect 16899 18921 16908 18955
rect 16856 18912 16908 18921
rect 7656 18708 7708 18760
rect 7932 18708 7984 18760
rect 9680 18708 9732 18760
rect 10140 18708 10192 18760
rect 10968 18751 11020 18760
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 4160 18640 4212 18692
rect 8668 18640 8720 18692
rect 1584 18615 1636 18624
rect 1584 18581 1593 18615
rect 1593 18581 1627 18615
rect 1627 18581 1636 18615
rect 1584 18572 1636 18581
rect 2136 18572 2188 18624
rect 8300 18572 8352 18624
rect 14924 18776 14976 18828
rect 12532 18708 12584 18760
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 14280 18751 14332 18760
rect 13268 18708 13320 18717
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 13452 18640 13504 18692
rect 15568 18708 15620 18760
rect 12900 18572 12952 18624
rect 14740 18572 14792 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 10600 18368 10652 18420
rect 14924 18411 14976 18420
rect 14924 18377 14933 18411
rect 14933 18377 14967 18411
rect 14967 18377 14976 18411
rect 14924 18368 14976 18377
rect 3516 18343 3568 18352
rect 3516 18309 3525 18343
rect 3525 18309 3559 18343
rect 3559 18309 3568 18343
rect 3516 18300 3568 18309
rect 4160 18300 4212 18352
rect 15292 18300 15344 18352
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 3240 18232 3292 18284
rect 7656 18232 7708 18284
rect 2688 18164 2740 18216
rect 7564 18164 7616 18216
rect 12808 18232 12860 18284
rect 14372 18232 14424 18284
rect 9772 18164 9824 18216
rect 2596 18028 2648 18080
rect 4988 18028 5040 18080
rect 10140 18028 10192 18080
rect 13452 18028 13504 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 4068 17688 4120 17740
rect 7748 17688 7800 17740
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 2136 17663 2188 17672
rect 2136 17629 2170 17663
rect 2170 17629 2188 17663
rect 2136 17620 2188 17629
rect 2412 17620 2464 17672
rect 7656 17620 7708 17672
rect 14832 17663 14884 17672
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3240 17484 3292 17493
rect 7380 17484 7432 17536
rect 7656 17484 7708 17536
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 16672 17663 16724 17672
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 14740 17595 14792 17604
rect 14740 17561 14749 17595
rect 14749 17561 14783 17595
rect 14783 17561 14792 17595
rect 14740 17552 14792 17561
rect 17224 17552 17276 17604
rect 15476 17484 15528 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 1400 17280 1452 17332
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 15292 17280 15344 17332
rect 16304 17280 16356 17332
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 9772 17187 9824 17196
rect 7380 17144 7432 17153
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 16672 17144 16724 17196
rect 16948 17144 17000 17196
rect 18144 17144 18196 17196
rect 11520 17076 11572 17128
rect 13636 17008 13688 17060
rect 7380 16940 7432 16992
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 12348 16940 12400 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7380 16779 7432 16788
rect 7380 16745 7389 16779
rect 7389 16745 7423 16779
rect 7423 16745 7432 16779
rect 7380 16736 7432 16745
rect 11520 16779 11572 16788
rect 11520 16745 11529 16779
rect 11529 16745 11563 16779
rect 11563 16745 11572 16779
rect 11520 16736 11572 16745
rect 16488 16779 16540 16788
rect 16488 16745 16497 16779
rect 16497 16745 16531 16779
rect 16531 16745 16540 16779
rect 16488 16736 16540 16745
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 1860 16600 1912 16652
rect 2780 16600 2832 16652
rect 2136 16532 2188 16584
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 5356 16464 5408 16516
rect 15476 16668 15528 16720
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 16304 16600 16356 16652
rect 9312 16532 9364 16584
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 10968 16532 11020 16584
rect 12348 16532 12400 16584
rect 16212 16532 16264 16584
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 2320 16396 2372 16448
rect 2504 16396 2556 16448
rect 7288 16396 7340 16448
rect 7840 16396 7892 16448
rect 10232 16464 10284 16516
rect 17776 16532 17828 16584
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 16672 16464 16724 16516
rect 17408 16396 17460 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 1676 16192 1728 16244
rect 2320 16167 2372 16176
rect 2320 16133 2354 16167
rect 2354 16133 2372 16167
rect 5356 16192 5408 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 17408 16192 17460 16201
rect 2320 16124 2372 16133
rect 1400 16056 1452 16108
rect 1860 16056 1912 16108
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 7656 16099 7708 16108
rect 6736 16056 6788 16065
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 8024 16056 8076 16108
rect 10232 16056 10284 16108
rect 13452 16124 13504 16176
rect 7288 15988 7340 16040
rect 5816 15920 5868 15972
rect 3424 15895 3476 15904
rect 3424 15861 3433 15895
rect 3433 15861 3467 15895
rect 3467 15861 3476 15895
rect 3424 15852 3476 15861
rect 5080 15852 5132 15904
rect 7380 15920 7432 15972
rect 11612 16056 11664 16108
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 16672 16056 16724 16108
rect 18052 16056 18104 16108
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11152 15852 11204 15904
rect 14648 15852 14700 15904
rect 16488 15852 16540 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 1492 15580 1544 15632
rect 6736 15580 6788 15632
rect 11612 15580 11664 15632
rect 14188 15648 14240 15700
rect 14648 15580 14700 15632
rect 15660 15648 15712 15700
rect 16488 15580 16540 15632
rect 2596 15555 2648 15564
rect 2596 15521 2605 15555
rect 2605 15521 2639 15555
rect 2639 15521 2648 15555
rect 2596 15512 2648 15521
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 7012 15512 7064 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 3424 15444 3476 15496
rect 7656 15487 7708 15496
rect 1860 15376 1912 15428
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 8208 15444 8260 15496
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 12164 15444 12216 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 16672 15444 16724 15496
rect 17316 15444 17368 15496
rect 17960 15444 18012 15496
rect 8300 15376 8352 15428
rect 1400 15351 1452 15360
rect 1400 15317 1409 15351
rect 1409 15317 1443 15351
rect 1443 15317 1452 15351
rect 1400 15308 1452 15317
rect 17868 15308 17920 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 17960 15104 18012 15156
rect 8300 15079 8352 15088
rect 8300 15045 8309 15079
rect 8309 15045 8343 15079
rect 8343 15045 8352 15079
rect 8300 15036 8352 15045
rect 1860 14968 1912 15020
rect 2320 14968 2372 15020
rect 7380 14968 7432 15020
rect 7564 14968 7616 15020
rect 10968 15036 11020 15088
rect 12256 14968 12308 15020
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 17500 15011 17552 15020
rect 17500 14977 17534 15011
rect 17534 14977 17552 15011
rect 17500 14968 17552 14977
rect 11244 14900 11296 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 17040 14900 17092 14952
rect 1584 14875 1636 14884
rect 1584 14841 1593 14875
rect 1593 14841 1627 14875
rect 1627 14841 1636 14875
rect 1584 14832 1636 14841
rect 1952 14832 2004 14884
rect 10324 14832 10376 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 9220 14764 9272 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14603 2372 14612
rect 2320 14569 2329 14603
rect 2329 14569 2363 14603
rect 2363 14569 2372 14603
rect 2320 14560 2372 14569
rect 2688 14560 2740 14612
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 10508 14560 10560 14612
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 16488 14560 16540 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 2596 14492 2648 14544
rect 1400 14424 1452 14476
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 5816 14467 5868 14476
rect 5816 14433 5825 14467
rect 5825 14433 5859 14467
rect 5859 14433 5868 14467
rect 5816 14424 5868 14433
rect 6276 14424 6328 14476
rect 15476 14424 15528 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 8760 14356 8812 14408
rect 9220 14399 9272 14408
rect 9220 14365 9254 14399
rect 9254 14365 9272 14399
rect 9220 14356 9272 14365
rect 10876 14399 10928 14408
rect 10876 14365 10885 14399
rect 10885 14365 10919 14399
rect 10919 14365 10928 14399
rect 10876 14356 10928 14365
rect 12900 14356 12952 14408
rect 14280 14356 14332 14408
rect 14464 14356 14516 14408
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 18236 14356 18288 14408
rect 2688 14263 2740 14272
rect 2688 14229 2697 14263
rect 2697 14229 2731 14263
rect 2731 14229 2740 14263
rect 2688 14220 2740 14229
rect 3976 14288 4028 14340
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 4620 14220 4672 14272
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 5724 14263 5776 14272
rect 5724 14229 5733 14263
rect 5733 14229 5767 14263
rect 5767 14229 5776 14263
rect 5724 14220 5776 14229
rect 13636 14220 13688 14272
rect 16856 14220 16908 14272
rect 17224 14220 17276 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2044 14016 2096 14068
rect 2228 13991 2280 14000
rect 2228 13957 2262 13991
rect 2262 13957 2280 13991
rect 2228 13948 2280 13957
rect 2688 14016 2740 14068
rect 8484 14016 8536 14068
rect 12716 14016 12768 14068
rect 13452 14016 13504 14068
rect 1768 13880 1820 13932
rect 3976 13880 4028 13932
rect 5356 13880 5408 13932
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 14096 13880 14148 13932
rect 2964 13812 3016 13864
rect 6276 13812 6328 13864
rect 9772 13812 9824 13864
rect 10232 13812 10284 13864
rect 10508 13812 10560 13864
rect 14280 13880 14332 13932
rect 16856 14016 16908 14068
rect 16948 13923 17000 13932
rect 16948 13889 16982 13923
rect 16982 13889 17000 13923
rect 16948 13880 17000 13889
rect 5816 13676 5868 13728
rect 13912 13676 13964 13728
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 16856 13676 16908 13728
rect 17040 13676 17092 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2412 13472 2464 13524
rect 5632 13472 5684 13524
rect 5724 13472 5776 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 10508 13472 10560 13524
rect 14096 13515 14148 13524
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 16948 13472 17000 13524
rect 3516 13268 3568 13320
rect 3976 13175 4028 13184
rect 3976 13141 3985 13175
rect 3985 13141 4019 13175
rect 4019 13141 4028 13175
rect 3976 13132 4028 13141
rect 5724 13311 5776 13320
rect 5724 13277 5747 13311
rect 5747 13277 5776 13311
rect 5724 13268 5776 13277
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 9680 13268 9732 13320
rect 10048 13268 10100 13320
rect 10508 13336 10560 13388
rect 13912 13336 13964 13388
rect 10876 13268 10928 13320
rect 12900 13268 12952 13320
rect 13176 13268 13228 13320
rect 13360 13268 13412 13320
rect 13728 13268 13780 13320
rect 15568 13268 15620 13320
rect 17224 13311 17276 13320
rect 5540 13132 5592 13184
rect 5632 13132 5684 13184
rect 9404 13132 9456 13184
rect 10508 13132 10560 13184
rect 15016 13200 15068 13252
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 17500 13268 17552 13320
rect 17132 13200 17184 13252
rect 15844 13132 15896 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 9404 12928 9456 12980
rect 15844 12928 15896 12980
rect 12348 12860 12400 12912
rect 14648 12903 14700 12912
rect 14648 12869 14657 12903
rect 14657 12869 14691 12903
rect 14691 12869 14700 12903
rect 14648 12860 14700 12869
rect 17132 12860 17184 12912
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 5724 12792 5776 12844
rect 6276 12724 6328 12776
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 4620 12588 4672 12640
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 7656 12792 7708 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 10140 12792 10192 12844
rect 6460 12724 6512 12776
rect 6552 12656 6604 12708
rect 7380 12588 7432 12640
rect 12900 12792 12952 12844
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 10324 12588 10376 12640
rect 13728 12656 13780 12708
rect 15292 12792 15344 12844
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 16948 12792 17000 12844
rect 16856 12724 16908 12776
rect 15384 12588 15436 12640
rect 17316 12588 17368 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2412 12384 2464 12436
rect 6460 12384 6512 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 12348 12384 12400 12436
rect 2596 12248 2648 12300
rect 13176 12384 13228 12436
rect 15384 12384 15436 12436
rect 16948 12427 17000 12436
rect 16948 12393 16957 12427
rect 16957 12393 16991 12427
rect 16991 12393 17000 12427
rect 16948 12384 17000 12393
rect 13268 12316 13320 12368
rect 13452 12316 13504 12368
rect 1400 12180 1452 12232
rect 4620 12180 4672 12232
rect 6092 12180 6144 12232
rect 8760 12180 8812 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 11704 12223 11756 12232
rect 11704 12189 11713 12223
rect 11713 12189 11747 12223
rect 11747 12189 11756 12223
rect 11704 12180 11756 12189
rect 3240 12112 3292 12164
rect 5632 12112 5684 12164
rect 12716 12180 12768 12232
rect 13360 12180 13412 12232
rect 15292 12180 15344 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 4344 12087 4396 12096
rect 2688 12044 2740 12053
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 16672 12112 16724 12164
rect 12532 12044 12584 12096
rect 13636 12044 13688 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 1860 11840 1912 11892
rect 2228 11772 2280 11824
rect 4344 11772 4396 11824
rect 1768 11704 1820 11756
rect 2504 11704 2556 11756
rect 5540 11704 5592 11756
rect 6092 11704 6144 11756
rect 12532 11840 12584 11892
rect 13636 11883 13688 11892
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 10324 11772 10376 11824
rect 7656 11704 7708 11756
rect 8668 11704 8720 11756
rect 9312 11704 9364 11756
rect 13360 11704 13412 11756
rect 14648 11772 14700 11824
rect 16764 11772 16816 11824
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 15936 11636 15988 11688
rect 6828 11568 6880 11620
rect 9772 11568 9824 11620
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 11244 11500 11296 11552
rect 11980 11500 12032 11552
rect 13360 11500 13412 11552
rect 18696 11568 18748 11620
rect 15384 11500 15436 11552
rect 17868 11500 17920 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13176 11296 13228 11348
rect 15936 11339 15988 11348
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 1584 11271 1636 11280
rect 1584 11237 1593 11271
rect 1593 11237 1627 11271
rect 1627 11237 1636 11271
rect 1584 11228 1636 11237
rect 3056 11228 3108 11280
rect 3240 11228 3292 11280
rect 11704 11228 11756 11280
rect 12532 11228 12584 11280
rect 2780 11092 2832 11144
rect 5816 11092 5868 11144
rect 8668 11092 8720 11144
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 12624 11135 12676 11144
rect 9312 11067 9364 11076
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 16856 11092 16908 11144
rect 10876 11024 10928 11076
rect 15292 11024 15344 11076
rect 17592 11067 17644 11076
rect 17592 11033 17626 11067
rect 17626 11033 17644 11067
rect 17592 11024 17644 11033
rect 12440 10956 12492 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 2688 10752 2740 10804
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 12808 10752 12860 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 15660 10795 15712 10804
rect 15660 10761 15669 10795
rect 15669 10761 15703 10795
rect 15703 10761 15712 10795
rect 15660 10752 15712 10761
rect 17592 10752 17644 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 1400 10616 1452 10668
rect 3884 10616 3936 10668
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 12072 10616 12124 10668
rect 17132 10684 17184 10736
rect 16580 10616 16632 10668
rect 19340 10616 19392 10668
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 11428 10548 11480 10600
rect 2872 10412 2924 10464
rect 9588 10412 9640 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 8668 10208 8720 10260
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 5632 10140 5684 10192
rect 5080 10072 5132 10124
rect 5356 10072 5408 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3332 10004 3384 10056
rect 5724 10004 5776 10056
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 8116 10047 8168 10056
rect 6092 10004 6144 10013
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 11980 10004 12032 10056
rect 14004 10004 14056 10056
rect 6368 9979 6420 9988
rect 6368 9945 6402 9979
rect 6402 9945 6420 9979
rect 6368 9936 6420 9945
rect 6552 9936 6604 9988
rect 2780 9868 2832 9920
rect 8852 9868 8904 9920
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 12440 9868 12492 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 2780 9639 2832 9648
rect 2780 9605 2814 9639
rect 2814 9605 2832 9639
rect 2780 9596 2832 9605
rect 6092 9528 6144 9580
rect 6184 9528 6236 9580
rect 8024 9528 8076 9580
rect 10048 9571 10100 9580
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 2504 9460 2556 9469
rect 7840 9460 7892 9512
rect 10048 9537 10057 9571
rect 10057 9537 10091 9571
rect 10091 9537 10100 9571
rect 10048 9528 10100 9537
rect 19248 9596 19300 9648
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16028 9528 16080 9580
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 8852 9435 8904 9444
rect 8852 9401 8861 9435
rect 8861 9401 8895 9435
rect 8895 9401 8904 9435
rect 8852 9392 8904 9401
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 5816 9324 5868 9376
rect 16488 9460 16540 9512
rect 11428 9392 11480 9444
rect 12532 9392 12584 9444
rect 16120 9324 16172 9376
rect 16856 9324 16908 9376
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9120 1728 9172
rect 5816 9120 5868 9172
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 2964 9052 3016 9104
rect 3240 9095 3292 9104
rect 3240 9061 3249 9095
rect 3249 9061 3283 9095
rect 3283 9061 3292 9095
rect 3240 9052 3292 9061
rect 5632 9095 5684 9104
rect 5632 9061 5641 9095
rect 5641 9061 5675 9095
rect 5675 9061 5684 9095
rect 5632 9052 5684 9061
rect 6092 9052 6144 9104
rect 10968 9120 11020 9172
rect 16028 9120 16080 9172
rect 19248 9163 19300 9172
rect 19248 9129 19257 9163
rect 19257 9129 19291 9163
rect 19291 9129 19300 9163
rect 19248 9120 19300 9129
rect 12256 9052 12308 9104
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2780 8916 2832 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3516 8916 3568 8968
rect 7748 8984 7800 9036
rect 10232 8984 10284 9036
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 8668 8916 8720 8968
rect 10048 8848 10100 8900
rect 11428 8916 11480 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 19156 8916 19208 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 20628 8916 20680 8968
rect 11520 8848 11572 8900
rect 12164 8848 12216 8900
rect 19064 8848 19116 8900
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 5908 8780 5960 8832
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19984 8780 20036 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 2044 8576 2096 8628
rect 11152 8576 11204 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11980 8576 12032 8628
rect 15568 8576 15620 8628
rect 15752 8576 15804 8628
rect 5724 8508 5776 8560
rect 6920 8508 6972 8560
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 8116 8551 8168 8560
rect 8116 8517 8125 8551
rect 8125 8517 8159 8551
rect 8159 8517 8168 8551
rect 8116 8508 8168 8517
rect 13176 8508 13228 8560
rect 19064 8576 19116 8628
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2504 8440 2556 8492
rect 5908 8440 5960 8492
rect 8668 8440 8720 8492
rect 10232 8440 10284 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 15936 8440 15988 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 18052 8508 18104 8560
rect 17316 8440 17368 8492
rect 18788 8508 18840 8560
rect 19984 8508 20036 8560
rect 19432 8440 19484 8492
rect 10508 8372 10560 8424
rect 11428 8372 11480 8424
rect 20444 8440 20496 8492
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 16212 8304 16264 8356
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4620 8236 4672 8288
rect 8116 8236 8168 8288
rect 8300 8236 8352 8288
rect 13084 8236 13136 8288
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1952 8032 2004 8084
rect 3976 8032 4028 8084
rect 7748 8032 7800 8084
rect 10508 8032 10560 8084
rect 11888 8032 11940 8084
rect 13360 8032 13412 8084
rect 8300 7964 8352 8016
rect 13084 7964 13136 8016
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3240 7896 3292 7948
rect 8208 7896 8260 7948
rect 6552 7828 6604 7880
rect 10324 7828 10376 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 3792 7692 3844 7744
rect 7104 7760 7156 7812
rect 8576 7760 8628 7812
rect 11152 7896 11204 7948
rect 16488 7896 16540 7948
rect 17868 7939 17920 7948
rect 17868 7905 17877 7939
rect 17877 7905 17911 7939
rect 17911 7905 17920 7939
rect 17868 7896 17920 7905
rect 17132 7828 17184 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 19984 7896 20036 7948
rect 20536 7828 20588 7880
rect 10600 7692 10652 7744
rect 13084 7692 13136 7744
rect 13820 7692 13872 7744
rect 14372 7692 14424 7744
rect 15016 7692 15068 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 3056 7488 3108 7540
rect 5908 7488 5960 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 7932 7488 7984 7540
rect 13820 7531 13872 7540
rect 2872 7420 2924 7472
rect 2412 7352 2464 7404
rect 4620 7420 4672 7472
rect 7472 7420 7524 7472
rect 3332 7352 3384 7404
rect 6000 7352 6052 7404
rect 6920 7395 6972 7404
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 3148 7284 3200 7336
rect 4804 7284 4856 7336
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7288 7352 7340 7404
rect 7840 7352 7892 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8852 7395 8904 7404
rect 8668 7352 8720 7361
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 5448 7216 5500 7268
rect 9772 7284 9824 7336
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 10784 7284 10836 7336
rect 13820 7497 13829 7531
rect 13829 7497 13863 7531
rect 13863 7497 13872 7531
rect 13820 7488 13872 7497
rect 14464 7488 14516 7540
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 13820 7352 13872 7404
rect 14648 7352 14700 7404
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 19248 7352 19300 7404
rect 13084 7284 13136 7336
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 6552 7148 6604 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 13820 7216 13872 7268
rect 14372 7148 14424 7200
rect 15752 7148 15804 7200
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2872 6987 2924 6996
rect 2872 6953 2881 6987
rect 2881 6953 2915 6987
rect 2915 6953 2924 6987
rect 2872 6944 2924 6953
rect 4068 6944 4120 6996
rect 6000 6944 6052 6996
rect 7840 6944 7892 6996
rect 1952 6808 2004 6860
rect 6736 6808 6788 6860
rect 7656 6876 7708 6928
rect 13176 6944 13228 6996
rect 18420 6876 18472 6928
rect 37280 6876 37332 6928
rect 8852 6808 8904 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3976 6740 4028 6792
rect 4620 6740 4672 6792
rect 5448 6740 5500 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 2412 6672 2464 6724
rect 3516 6672 3568 6724
rect 2780 6604 2832 6656
rect 4804 6604 4856 6656
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7288 6740 7340 6792
rect 7656 6740 7708 6792
rect 14464 6808 14516 6860
rect 15752 6808 15804 6860
rect 17132 6851 17184 6860
rect 17132 6817 17141 6851
rect 17141 6817 17175 6851
rect 17175 6817 17184 6851
rect 17132 6808 17184 6817
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 15936 6740 15988 6792
rect 10416 6672 10468 6724
rect 16212 6740 16264 6792
rect 16304 6672 16356 6724
rect 10508 6604 10560 6656
rect 10600 6604 10652 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 10876 6400 10928 6452
rect 14556 6400 14608 6452
rect 15292 6400 15344 6452
rect 3332 6375 3384 6384
rect 3332 6341 3341 6375
rect 3341 6341 3375 6375
rect 3375 6341 3384 6375
rect 3332 6332 3384 6341
rect 6000 6332 6052 6384
rect 7380 6332 7432 6384
rect 2780 6264 2832 6316
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 11336 6332 11388 6384
rect 11704 6332 11756 6384
rect 13452 6332 13504 6384
rect 10876 6307 10928 6316
rect 3240 6196 3292 6248
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 13820 6264 13872 6316
rect 15660 6332 15712 6384
rect 16212 6332 16264 6384
rect 7196 6196 7248 6248
rect 16028 6264 16080 6316
rect 16396 6264 16448 6316
rect 38568 6264 38620 6316
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 5264 6128 5316 6180
rect 10692 6128 10744 6180
rect 16856 6128 16908 6180
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3976 5856 4028 5908
rect 9956 5856 10008 5908
rect 15200 5856 15252 5908
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 3240 5720 3292 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 16488 5788 16540 5840
rect 1492 5652 1544 5704
rect 1676 5652 1728 5704
rect 6828 5695 6880 5704
rect 6828 5661 6862 5695
rect 6862 5661 6880 5695
rect 6828 5652 6880 5661
rect 2596 5516 2648 5568
rect 3608 5516 3660 5568
rect 6184 5516 6236 5568
rect 6736 5516 6788 5568
rect 15016 5652 15068 5704
rect 15384 5652 15436 5704
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 15292 5584 15344 5636
rect 15384 5516 15436 5568
rect 16764 5559 16816 5568
rect 16764 5525 16773 5559
rect 16773 5525 16807 5559
rect 16807 5525 16816 5559
rect 16764 5516 16816 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 10692 5312 10744 5364
rect 13544 5312 13596 5364
rect 15108 5312 15160 5364
rect 15844 5312 15896 5364
rect 17776 5312 17828 5364
rect 6828 5244 6880 5296
rect 15292 5244 15344 5296
rect 16764 5244 16816 5296
rect 18880 5244 18932 5296
rect 19340 5244 19392 5296
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2320 5176 2372 5228
rect 2504 5219 2556 5228
rect 2504 5185 2538 5219
rect 2538 5185 2556 5219
rect 2504 5176 2556 5185
rect 4620 5176 4672 5228
rect 5448 5176 5500 5228
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 11152 5176 11204 5228
rect 3792 5108 3844 5160
rect 9864 5151 9916 5160
rect 3884 5040 3936 5092
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 10048 5108 10100 5160
rect 15108 5176 15160 5228
rect 15384 5219 15436 5228
rect 15384 5185 15393 5219
rect 15393 5185 15427 5219
rect 15427 5185 15436 5219
rect 15384 5176 15436 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 16856 5219 16908 5228
rect 15660 5176 15712 5185
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 30288 5176 30340 5228
rect 5724 4972 5776 5024
rect 8208 4972 8260 5024
rect 10508 5040 10560 5092
rect 10140 5015 10192 5024
rect 10140 4981 10149 5015
rect 10149 4981 10183 5015
rect 10183 4981 10192 5015
rect 10140 4972 10192 4981
rect 11520 4972 11572 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2504 4768 2556 4820
rect 9864 4768 9916 4820
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 14832 4768 14884 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 5448 4700 5500 4752
rect 3608 4632 3660 4684
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 3148 4564 3200 4616
rect 4160 4564 4212 4616
rect 5172 4564 5224 4616
rect 6552 4632 6604 4684
rect 5356 4496 5408 4548
rect 10048 4564 10100 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 16856 4632 16908 4684
rect 11612 4564 11664 4573
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 18788 4632 18840 4684
rect 18880 4632 18932 4684
rect 19064 4564 19116 4616
rect 24584 4607 24636 4616
rect 9772 4496 9824 4548
rect 16764 4496 16816 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4344 4428 4396 4480
rect 10232 4428 10284 4480
rect 18512 4428 18564 4480
rect 19340 4496 19392 4548
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 24676 4428 24728 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 10232 4224 10284 4276
rect 24584 4224 24636 4276
rect 7932 4156 7984 4208
rect 18512 4156 18564 4208
rect 2320 4088 2372 4140
rect 3148 4088 3200 4140
rect 3240 4088 3292 4140
rect 2688 4020 2740 4072
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 4344 4131 4396 4140
rect 3700 4088 3752 4097
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 3976 4020 4028 4072
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 9772 4131 9824 4140
rect 6828 4088 6880 4097
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 10232 4131 10284 4140
rect 3608 3952 3660 4004
rect 5264 3952 5316 4004
rect 204 3884 256 3936
rect 3884 3884 3936 3936
rect 4712 3884 4764 3936
rect 5080 3884 5132 3936
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 11244 4088 11296 4140
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 11336 4020 11388 4072
rect 16304 4020 16356 4072
rect 17592 4020 17644 4072
rect 19432 4088 19484 4140
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 25596 4088 25648 4140
rect 28816 4020 28868 4072
rect 10968 3952 11020 4004
rect 21272 3952 21324 4004
rect 6460 3884 6512 3936
rect 8392 3884 8444 3936
rect 11888 3884 11940 3936
rect 14832 3884 14884 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 664 3612 716 3664
rect 4804 3680 4856 3732
rect 9588 3680 9640 3732
rect 11612 3680 11664 3732
rect 16580 3723 16632 3732
rect 16580 3689 16589 3723
rect 16589 3689 16623 3723
rect 16623 3689 16632 3723
rect 16580 3680 16632 3689
rect 17500 3680 17552 3732
rect 15752 3612 15804 3664
rect 16120 3612 16172 3664
rect 3148 3544 3200 3596
rect 10784 3544 10836 3596
rect 3056 3476 3108 3528
rect 3884 3476 3936 3528
rect 6460 3519 6512 3528
rect 3700 3408 3752 3460
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 7472 3476 7524 3528
rect 10416 3476 10468 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 1584 3340 1636 3392
rect 2688 3340 2740 3392
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 6276 3340 6328 3349
rect 6368 3340 6420 3392
rect 10968 3340 11020 3392
rect 16304 3544 16356 3596
rect 12348 3476 12400 3528
rect 13360 3476 13412 3528
rect 14740 3476 14792 3528
rect 16212 3476 16264 3528
rect 16948 3544 17000 3596
rect 17592 3544 17644 3596
rect 18328 3476 18380 3528
rect 19708 3544 19760 3596
rect 18512 3476 18564 3528
rect 25688 3476 25740 3528
rect 11888 3408 11940 3460
rect 15200 3408 15252 3460
rect 59636 3408 59688 3460
rect 12624 3340 12676 3392
rect 12716 3340 12768 3392
rect 14924 3340 14976 3392
rect 16672 3340 16724 3392
rect 17040 3340 17092 3392
rect 17132 3340 17184 3392
rect 19984 3340 20036 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 2136 3136 2188 3188
rect 4068 3136 4120 3188
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 1952 3000 2004 3052
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 6184 3068 6236 3120
rect 6276 3068 6328 3120
rect 4620 3000 4672 3052
rect 5724 3043 5776 3052
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 2412 2932 2464 2984
rect 5080 2932 5132 2984
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 8208 3000 8260 3052
rect 6368 2932 6420 2984
rect 10876 3136 10928 3188
rect 11980 3136 12032 3188
rect 14004 3136 14056 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 18328 3136 18380 3188
rect 12624 3111 12676 3120
rect 9312 3000 9364 3052
rect 10600 3000 10652 3052
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 10784 3000 10836 3052
rect 10968 3043 11020 3052
rect 10968 3009 10977 3043
rect 10977 3009 11011 3043
rect 11011 3009 11020 3043
rect 10968 3000 11020 3009
rect 11428 3000 11480 3052
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 15752 3068 15804 3120
rect 12716 3000 12768 3009
rect 2596 2864 2648 2916
rect 3700 2864 3752 2916
rect 5632 2864 5684 2916
rect 11980 2864 12032 2916
rect 1124 2796 1176 2848
rect 1676 2796 1728 2848
rect 2872 2839 2924 2848
rect 2872 2805 2881 2839
rect 2881 2805 2915 2839
rect 2915 2805 2924 2839
rect 2872 2796 2924 2805
rect 3516 2796 3568 2848
rect 6368 2796 6420 2848
rect 9036 2796 9088 2848
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 11336 2796 11388 2848
rect 14740 3000 14792 3052
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15200 3000 15252 3052
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 17040 2932 17092 2984
rect 18972 3000 19024 3052
rect 19156 3068 19208 3120
rect 21272 3043 21324 3052
rect 18696 2932 18748 2984
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 23572 3000 23624 3052
rect 19984 2932 20036 2984
rect 56692 3000 56744 3052
rect 33324 2932 33376 2984
rect 17684 2864 17736 2916
rect 17960 2864 18012 2916
rect 22192 2864 22244 2916
rect 16672 2796 16724 2848
rect 16856 2796 16908 2848
rect 19432 2796 19484 2848
rect 20168 2796 20220 2848
rect 21640 2796 21692 2848
rect 25044 2796 25096 2848
rect 32312 2796 32364 2848
rect 35348 2796 35400 2848
rect 36728 2796 36780 2848
rect 39672 2796 39724 2848
rect 42616 2796 42668 2848
rect 44088 2796 44140 2848
rect 46940 2796 46992 2848
rect 49884 2796 49936 2848
rect 52828 2796 52880 2848
rect 54300 2796 54352 2848
rect 58716 2796 58768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10232 2592 10284 2644
rect 14372 2592 14424 2644
rect 5632 2524 5684 2576
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 6460 2456 6512 2508
rect 1308 2388 1360 2440
rect 4712 2388 4764 2440
rect 5540 2388 5592 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 8484 2388 8536 2440
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 17592 2524 17644 2576
rect 15292 2456 15344 2508
rect 16764 2499 16816 2508
rect 16764 2465 16773 2499
rect 16773 2465 16807 2499
rect 16807 2465 16816 2499
rect 16764 2456 16816 2465
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 14280 2388 14332 2440
rect 14832 2388 14884 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17960 2456 18012 2508
rect 19064 2592 19116 2644
rect 25596 2635 25648 2644
rect 18972 2524 19024 2576
rect 21180 2524 21232 2576
rect 25320 2524 25372 2576
rect 25596 2601 25605 2635
rect 25605 2601 25639 2635
rect 25639 2601 25648 2635
rect 25596 2592 25648 2601
rect 25688 2592 25740 2644
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 30288 2635 30340 2644
rect 30288 2601 30297 2635
rect 30297 2601 30331 2635
rect 30331 2601 30340 2635
rect 30288 2592 30340 2601
rect 37280 2592 37332 2644
rect 30472 2524 30524 2576
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 19156 2388 19208 2440
rect 19432 2388 19484 2440
rect 21088 2388 21140 2440
rect 21456 2456 21508 2508
rect 21548 2388 21600 2440
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22560 2388 22612 2440
rect 24032 2388 24084 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 25964 2388 26016 2440
rect 26516 2388 26568 2440
rect 27436 2388 27488 2440
rect 27988 2388 28040 2440
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30380 2388 30432 2440
rect 30840 2388 30892 2440
rect 31852 2388 31904 2440
rect 33784 2388 33836 2440
rect 34796 2388 34848 2440
rect 35164 2431 35216 2440
rect 35164 2397 35173 2431
rect 35173 2397 35207 2431
rect 35207 2397 35216 2431
rect 35164 2388 35216 2397
rect 15936 2320 15988 2372
rect 21180 2320 21232 2372
rect 38200 2388 38252 2440
rect 3056 2252 3108 2304
rect 6000 2252 6052 2304
rect 7932 2252 7984 2304
rect 8944 2252 8996 2304
rect 10876 2252 10928 2304
rect 11888 2252 11940 2304
rect 13820 2252 13872 2304
rect 14832 2252 14884 2304
rect 17224 2252 17276 2304
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 20076 2252 20128 2304
rect 36268 2320 36320 2372
rect 37740 2320 37792 2372
rect 38568 2320 38620 2372
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 41328 2388 41380 2440
rect 22100 2252 22152 2304
rect 24584 2252 24636 2304
rect 25320 2252 25372 2304
rect 40408 2295 40460 2304
rect 40408 2261 40417 2295
rect 40417 2261 40451 2295
rect 40451 2261 40460 2295
rect 40408 2252 40460 2261
rect 40500 2252 40552 2304
rect 42064 2320 42116 2372
rect 43076 2431 43128 2440
rect 43076 2397 43085 2431
rect 43085 2397 43119 2431
rect 43119 2397 43128 2431
rect 43076 2388 43128 2397
rect 43536 2388 43588 2440
rect 45008 2388 45060 2440
rect 45468 2388 45520 2440
rect 46480 2388 46532 2440
rect 47952 2388 48004 2440
rect 48412 2388 48464 2440
rect 49424 2388 49476 2440
rect 50896 2388 50948 2440
rect 51356 2388 51408 2440
rect 52368 2388 52420 2440
rect 53840 2388 53892 2440
rect 55220 2388 55272 2440
rect 55772 2388 55824 2440
rect 57244 2388 57296 2440
rect 46756 2295 46808 2304
rect 46756 2261 46765 2295
rect 46765 2261 46799 2295
rect 46799 2261 46808 2295
rect 46756 2252 46808 2261
rect 58164 2320 58216 2372
rect 48320 2252 48372 2304
rect 51172 2295 51224 2304
rect 51172 2261 51181 2295
rect 51181 2261 51215 2295
rect 51215 2261 51224 2295
rect 51172 2252 51224 2261
rect 52920 2295 52972 2304
rect 52920 2261 52929 2295
rect 52929 2261 52963 2295
rect 52963 2261 52972 2295
rect 52920 2252 52972 2261
rect 55496 2295 55548 2304
rect 55496 2261 55505 2295
rect 55505 2261 55539 2295
rect 55539 2261 55548 2295
rect 55496 2252 55548 2261
rect 57060 2295 57112 2304
rect 57060 2261 57069 2295
rect 57069 2261 57103 2295
rect 57103 2261 57112 2295
rect 57060 2252 57112 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 14556 2048 14608 2100
rect 21456 2048 21508 2100
rect 21548 2048 21600 2100
rect 46756 2048 46808 2100
rect 15660 1980 15712 2032
rect 20076 1980 20128 2032
rect 20812 1980 20864 2032
rect 51172 1980 51224 2032
rect 15016 1912 15068 1964
rect 43076 1912 43128 1964
rect 15108 1844 15160 1896
rect 40408 1844 40460 1896
rect 20628 1776 20680 1828
rect 30472 1776 30524 1828
rect 17316 1708 17368 1760
rect 57060 1708 57112 1760
rect 20536 1640 20588 1692
rect 55496 1640 55548 1692
rect 15844 1572 15896 1624
rect 35164 1572 35216 1624
rect 20444 1504 20496 1556
rect 52920 1504 52972 1556
rect 2780 1436 2832 1488
rect 5172 1436 5224 1488
rect 19248 1436 19300 1488
rect 48320 1436 48372 1488
rect 16028 1368 16080 1420
rect 40500 1368 40552 1420
rect 3424 1164 3476 1216
rect 7104 1164 7156 1216
<< metal2 >>
rect 2778 41712 2834 41721
rect 2778 41647 2834 41656
rect 1582 40896 1638 40905
rect 1582 40831 1638 40840
rect 1490 40080 1546 40089
rect 1490 40015 1546 40024
rect 1504 38554 1532 40015
rect 1596 39642 1624 40831
rect 2792 39642 2820 41647
rect 3698 41200 3754 42000
rect 11150 41200 11206 42000
rect 18694 41200 18750 42000
rect 26146 41200 26202 42000
rect 33690 41200 33746 42000
rect 41142 41200 41198 42000
rect 48686 41200 48742 42000
rect 56138 41200 56194 42000
rect 3712 39642 3740 41200
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 1584 39636 1636 39642
rect 1584 39578 1636 39584
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 3700 39636 3752 39642
rect 3700 39578 3752 39584
rect 18708 39506 18736 41200
rect 26160 39658 26188 41200
rect 41156 39930 41184 41200
rect 41156 39902 41460 39930
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 26160 39642 26280 39658
rect 41432 39642 41460 39902
rect 48700 39642 48728 41200
rect 56152 39642 56180 41200
rect 26160 39636 26292 39642
rect 26160 39630 26240 39636
rect 26240 39578 26292 39584
rect 41420 39636 41472 39642
rect 41420 39578 41472 39584
rect 48688 39636 48740 39642
rect 48688 39578 48740 39584
rect 56140 39636 56192 39642
rect 56140 39578 56192 39584
rect 18696 39500 18748 39506
rect 18696 39442 18748 39448
rect 2136 39432 2188 39438
rect 2136 39374 2188 39380
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 1584 38752 1636 38758
rect 1584 38694 1636 38700
rect 1492 38548 1544 38554
rect 1492 38490 1544 38496
rect 1596 38457 1624 38694
rect 1582 38448 1638 38457
rect 1582 38383 1638 38392
rect 1492 38344 1544 38350
rect 1492 38286 1544 38292
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 26625 1440 28018
rect 1398 26616 1454 26625
rect 1398 26551 1454 26560
rect 1400 24064 1452 24070
rect 1400 24006 1452 24012
rect 1412 21706 1440 24006
rect 1504 22778 1532 38286
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 1584 37664 1636 37670
rect 1582 37632 1584 37641
rect 1636 37632 1638 37641
rect 1582 37567 1638 37576
rect 1582 36680 1638 36689
rect 1582 36615 1584 36624
rect 1636 36615 1638 36624
rect 1584 36586 1636 36592
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35873 1624 35974
rect 1582 35864 1638 35873
rect 1582 35799 1638 35808
rect 1582 35048 1638 35057
rect 1582 34983 1638 34992
rect 1596 34950 1624 34983
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 34241 1624 34546
rect 1582 34232 1638 34241
rect 1582 34167 1638 34176
rect 1584 33856 1636 33862
rect 1582 33824 1584 33833
rect 1636 33824 1638 33833
rect 1582 33759 1638 33768
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1596 33017 1624 33458
rect 1582 33008 1638 33017
rect 1582 32943 1638 32952
rect 1584 32564 1636 32570
rect 1584 32506 1636 32512
rect 1596 32473 1624 32506
rect 1582 32464 1638 32473
rect 1582 32399 1638 32408
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 1596 31657 1624 31758
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1582 31240 1638 31249
rect 1582 31175 1584 31184
rect 1636 31175 1638 31184
rect 1584 31146 1636 31152
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 1596 30433 1624 30670
rect 1582 30424 1638 30433
rect 1582 30359 1638 30368
rect 1584 30048 1636 30054
rect 1582 30016 1584 30025
rect 1636 30016 1638 30025
rect 1582 29951 1638 29960
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 1596 29209 1624 29582
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1584 29028 1636 29034
rect 1584 28970 1636 28976
rect 1596 28801 1624 28970
rect 1582 28792 1638 28801
rect 1582 28727 1638 28736
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1596 27334 1624 27367
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1584 26240 1636 26246
rect 1582 26208 1584 26217
rect 1636 26208 1638 26217
rect 1582 26143 1638 26152
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1596 25401 1624 25842
rect 1582 25392 1638 25401
rect 1582 25327 1638 25336
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 24993 1624 25094
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24177 1624 24754
rect 1582 24168 1638 24177
rect 1582 24103 1638 24112
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1596 23769 1624 23802
rect 1582 23760 1638 23769
rect 1582 23695 1638 23704
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1596 22817 1624 23054
rect 1582 22808 1638 22817
rect 1492 22772 1544 22778
rect 1582 22743 1638 22752
rect 1492 22714 1544 22720
rect 1492 22636 1544 22642
rect 1492 22578 1544 22584
rect 1320 21678 1440 21706
rect 1320 19258 1348 21678
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 1412 20942 1440 21519
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1398 20360 1454 20369
rect 1398 20295 1454 20304
rect 1412 19378 1440 20295
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1320 19230 1440 19258
rect 1412 17338 1440 19230
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 1412 16114 1440 16487
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1504 15638 1532 22578
rect 1584 22432 1636 22438
rect 1582 22400 1584 22409
rect 1636 22400 1638 22409
rect 1582 22335 1638 22344
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 21185 1624 21286
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1584 19984 1636 19990
rect 1582 19952 1584 19961
rect 1636 19952 1638 19961
rect 1582 19887 1638 19896
rect 1584 18624 1636 18630
rect 1582 18592 1584 18601
rect 1636 18592 1638 18601
rect 1582 18527 1638 18536
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17785 1624 18226
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1582 17368 1638 17377
rect 1582 17303 1584 17312
rect 1636 17303 1638 17312
rect 1584 17274 1636 17280
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16153 1624 16390
rect 1688 16250 1716 37810
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1780 24070 1808 36722
rect 1860 36168 1912 36174
rect 1860 36110 1912 36116
rect 1872 24070 1900 36110
rect 2148 35894 2176 39374
rect 2320 39364 2372 39370
rect 2320 39306 2372 39312
rect 2056 35866 2176 35894
rect 1952 35080 2004 35086
rect 1952 35022 2004 35028
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1964 23882 1992 35022
rect 1780 23854 1992 23882
rect 1780 18834 1808 23854
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 18970 1900 23666
rect 1952 22772 2004 22778
rect 1952 22714 2004 22720
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1872 16658 1900 17614
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1582 16144 1638 16153
rect 1872 16114 1900 16594
rect 1582 16079 1638 16088
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1492 15632 1544 15638
rect 1492 15574 1544 15580
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1400 15360 1452 15366
rect 1596 15337 1624 15438
rect 1872 15434 1900 16050
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1400 15302 1452 15308
rect 1582 15328 1638 15337
rect 1412 14482 1440 15302
rect 1582 15263 1638 15272
rect 1872 15178 1900 15370
rect 1780 15150 1900 15178
rect 1582 14920 1638 14929
rect 1582 14855 1584 14864
rect 1636 14855 1638 14864
rect 1584 14826 1636 14832
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1596 13977 1624 14350
rect 1582 13968 1638 13977
rect 1780 13938 1808 15150
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1582 13903 1638 13912
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1582 13560 1638 13569
rect 1582 13495 1584 13504
rect 1636 13495 1638 13504
rect 1584 13466 1636 13472
rect 1398 12744 1454 12753
rect 1398 12679 1454 12688
rect 1412 12238 1440 12679
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1780 11762 1808 13874
rect 1872 11898 1900 14962
rect 1964 14890 1992 22714
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 2056 14074 2084 35866
rect 2136 33312 2188 33318
rect 2136 33254 2188 33260
rect 2148 32910 2176 33254
rect 2136 32904 2188 32910
rect 2136 32846 2188 32852
rect 2332 28642 2360 39306
rect 3056 39296 3108 39302
rect 3054 39264 3056 39273
rect 3108 39264 3110 39273
rect 3054 39199 3110 39208
rect 2504 38956 2556 38962
rect 2504 38898 2556 38904
rect 2516 35894 2544 38898
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 6656 35894 6684 39374
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 2516 35866 2636 35894
rect 6656 35866 6776 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 2412 33516 2464 33522
rect 2412 33458 2464 33464
rect 2424 32570 2452 33458
rect 2412 32564 2464 32570
rect 2412 32506 2464 32512
rect 2504 28960 2556 28966
rect 2504 28902 2556 28908
rect 2332 28614 2452 28642
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2332 28218 2360 28426
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2228 27328 2280 27334
rect 2228 27270 2280 27276
rect 2240 27062 2268 27270
rect 2228 27056 2280 27062
rect 2228 26998 2280 27004
rect 2332 26586 2360 27406
rect 2320 26580 2372 26586
rect 2320 26522 2372 26528
rect 2424 26234 2452 28614
rect 2516 28082 2544 28902
rect 2608 28082 2636 35866
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 2872 34740 2924 34746
rect 2872 34682 2924 34688
rect 2780 32836 2832 32842
rect 2780 32778 2832 32784
rect 2792 32298 2820 32778
rect 2884 32570 2912 34682
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 4988 33380 5040 33386
rect 4988 33322 5040 33328
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 4632 32502 4660 32982
rect 5000 32978 5028 33322
rect 4988 32972 5040 32978
rect 4988 32914 5040 32920
rect 5080 32972 5132 32978
rect 5080 32914 5132 32920
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4620 32496 4672 32502
rect 4620 32438 4672 32444
rect 3148 32360 3200 32366
rect 3148 32302 3200 32308
rect 2780 32292 2832 32298
rect 2780 32234 2832 32240
rect 2792 31278 2820 32234
rect 2964 31952 3016 31958
rect 2964 31894 3016 31900
rect 2872 31680 2924 31686
rect 2872 31622 2924 31628
rect 2884 31414 2912 31622
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29850 2728 30194
rect 2792 30122 2820 31214
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 2884 30734 2912 31078
rect 2976 30802 3004 31894
rect 3056 31816 3108 31822
rect 3056 31758 3108 31764
rect 3068 30938 3096 31758
rect 3056 30932 3108 30938
rect 3056 30874 3108 30880
rect 3160 30802 3188 32302
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 31414 4660 32438
rect 4712 32428 4764 32434
rect 4712 32370 4764 32376
rect 4724 32026 4752 32370
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 4816 31822 4844 32710
rect 4908 32570 4936 32710
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4804 31816 4856 31822
rect 4804 31758 4856 31764
rect 4620 31408 4672 31414
rect 4620 31350 4672 31356
rect 4908 31346 4936 32506
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4988 31340 5040 31346
rect 4988 31282 5040 31288
rect 2964 30796 3016 30802
rect 2964 30738 3016 30744
rect 3148 30796 3200 30802
rect 3148 30738 3200 30744
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2780 30116 2832 30122
rect 2780 30058 2832 30064
rect 2964 30116 3016 30122
rect 2964 30058 3016 30064
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 2884 29306 2912 29446
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2780 29164 2832 29170
rect 2780 29106 2832 29112
rect 2688 29096 2740 29102
rect 2688 29038 2740 29044
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2700 28014 2728 29038
rect 2792 28422 2820 29106
rect 2976 28558 3004 30058
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2780 28416 2832 28422
rect 2780 28358 2832 28364
rect 2688 28008 2740 28014
rect 2608 27956 2688 27962
rect 2608 27950 2740 27956
rect 2504 27940 2556 27946
rect 2504 27882 2556 27888
rect 2608 27934 2728 27950
rect 2332 26206 2452 26234
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 24206 2176 24550
rect 2136 24200 2188 24206
rect 2136 24142 2188 24148
rect 2136 24064 2188 24070
rect 2136 24006 2188 24012
rect 2148 23746 2176 24006
rect 2240 23866 2268 24754
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2148 23718 2268 23746
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2148 22030 2176 22374
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2240 21842 2268 23718
rect 2148 21814 2268 21842
rect 2148 19922 2176 21814
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20534 2268 20742
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2240 19145 2268 19314
rect 2226 19136 2282 19145
rect 2226 19071 2282 19080
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 17678 2176 18566
rect 2240 18426 2268 18702
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2136 16584 2188 16590
rect 2332 16574 2360 26206
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2424 21690 2452 22578
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2424 20058 2452 20878
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2424 17678 2452 19858
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2332 16546 2452 16574
rect 2136 16526 2188 16532
rect 2148 15706 2176 16526
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16182 2360 16390
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2240 14006 2268 14758
rect 2332 14618 2360 14962
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2424 13530 2452 16546
rect 2516 16454 2544 27882
rect 2608 26330 2636 27934
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2700 26450 2728 27814
rect 2976 27402 3004 28494
rect 3054 27840 3110 27849
rect 3054 27775 3110 27784
rect 3068 27470 3096 27775
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 2964 27396 3016 27402
rect 2964 27338 3016 27344
rect 2976 26994 3004 27338
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 3160 26586 3188 26726
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2872 26444 2924 26450
rect 2872 26386 2924 26392
rect 2884 26330 2912 26386
rect 2608 26302 2912 26330
rect 3160 26314 3188 26522
rect 3148 26308 3200 26314
rect 2608 24750 2636 26302
rect 3148 26250 3200 26256
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2608 23746 2636 24686
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2700 23866 2728 24618
rect 2792 24138 2820 25230
rect 2780 24132 2832 24138
rect 2780 24074 2832 24080
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2608 23718 2728 23746
rect 2700 23662 2728 23718
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2792 23118 2820 24074
rect 3332 24064 3384 24070
rect 3332 24006 3384 24012
rect 3344 23730 3372 24006
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2608 21418 2636 22510
rect 2792 21962 2820 23054
rect 2780 21956 2832 21962
rect 2780 21898 2832 21904
rect 2688 21480 2740 21486
rect 2688 21422 2740 21428
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2608 19922 2636 21354
rect 2700 21146 2728 21422
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2792 20466 2820 21898
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21554 3280 21830
rect 3344 21554 3372 23666
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2608 18306 2636 19858
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2700 19514 2728 19654
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2792 19378 2820 20402
rect 3344 19786 3372 20538
rect 3332 19780 3384 19786
rect 3332 19722 3384 19728
rect 3436 19514 3464 31282
rect 4620 31204 4672 31210
rect 4620 31146 4672 31152
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3620 24818 3648 25638
rect 3712 25294 3740 27406
rect 3804 26314 3832 28358
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3896 27334 3924 28018
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3988 27674 4016 27950
rect 4068 27872 4120 27878
rect 4068 27814 4120 27820
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4080 27554 4108 27814
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4080 27526 4200 27554
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 3896 26450 3924 27270
rect 3988 27130 4016 27338
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 4172 26994 4200 27526
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 3792 26308 3844 26314
rect 3792 26250 3844 26256
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3700 25288 3752 25294
rect 3700 25230 3752 25236
rect 3896 24954 3924 25842
rect 3988 25498 4016 26318
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 3988 24886 4016 25434
rect 4080 25226 4108 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 3976 24880 4028 24886
rect 3976 24822 4028 24828
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18426 2728 19110
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2608 18278 2728 18306
rect 2700 18222 2728 18278
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2608 15570 2636 18022
rect 2700 15570 2728 18158
rect 2792 16658 2820 19314
rect 3528 18358 3556 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23202 4660 31146
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4724 29578 4752 30534
rect 4908 29714 4936 30738
rect 5000 30394 5028 31282
rect 5092 30802 5120 32914
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 4896 29708 4948 29714
rect 4896 29650 4948 29656
rect 4712 29572 4764 29578
rect 4712 29514 4764 29520
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 4724 24154 4752 26454
rect 4724 24126 4844 24154
rect 4632 23174 4752 23202
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3896 22778 3924 22918
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 3988 22710 4016 22918
rect 3700 22704 3752 22710
rect 3700 22646 3752 22652
rect 3976 22704 4028 22710
rect 3976 22646 4028 22652
rect 3712 21554 3740 22646
rect 4080 22166 4108 23054
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22778 4660 22986
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 4724 22098 4752 23174
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21690 4016 21966
rect 4816 21962 4844 24126
rect 4908 22094 4936 29650
rect 5000 29646 5028 30330
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 4908 22066 5028 22094
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3804 20602 3832 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4724 21010 4752 21830
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4080 18766 4108 19314
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 17542 3280 18226
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2700 14618 2728 15506
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 2240 11830 2268 12582
rect 2424 12442 2452 12786
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2608 12306 2636 14486
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 14074 2728 14214
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2976 13870 3004 14418
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3252 12434 3280 17478
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3436 15502 3464 15846
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3528 13326 3556 18294
rect 4080 17746 4108 18702
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4172 18358 4200 18634
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 3988 13938 4016 14282
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3252 12406 3372 12434
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 3240 12164 3292 12170
rect 3240 12106 3292 12112
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 1398 11520 1454 11529
rect 1398 11455 1454 11464
rect 1412 10674 1440 11455
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1596 11121 1624 11222
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1412 9897 1440 9998
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1688 9178 1716 9998
rect 2516 9518 2544 11698
rect 2700 10810 2728 12038
rect 3252 11558 3280 12106
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11286 3280 11494
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2792 10305 2820 11086
rect 3068 10810 3096 11222
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2884 10062 2912 10406
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9654 2820 9862
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8537 1624 8910
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 8634 2084 8774
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1582 8528 1638 8537
rect 2516 8498 2544 9454
rect 3252 9110 3280 10542
rect 3344 10062 3372 12406
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 1582 8463 1638 8472
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1964 8090 1992 8434
rect 2792 8129 2820 8910
rect 2778 8120 2834 8129
rect 1952 8084 2004 8090
rect 2778 8055 2834 8064
rect 1952 8026 2004 8032
rect 2976 7954 3004 9046
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 1584 7744 1636 7750
rect 1582 7712 1584 7721
rect 1636 7712 1638 7721
rect 1582 7647 1638 7656
rect 3068 7546 3096 8910
rect 3252 7954 3280 9046
rect 3528 8974 3556 13262
rect 3988 13190 4016 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 9382 3924 10610
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1490 6896 1546 6905
rect 1964 6866 1992 7278
rect 1490 6831 1546 6840
rect 1952 6860 2004 6866
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6497 1440 6734
rect 1398 6488 1454 6497
rect 1398 6423 1454 6432
rect 1504 5710 1532 6831
rect 1952 6802 2004 6808
rect 1584 6112 1636 6118
rect 1582 6080 1584 6089
rect 1636 6080 1638 6089
rect 1582 6015 1638 6024
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4729 1624 5170
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4321 1624 4422
rect 1582 4312 1638 4321
rect 1582 4247 1638 4256
rect 204 3936 256 3942
rect 204 3878 256 3884
rect 216 800 244 3878
rect 664 3664 716 3670
rect 664 3606 716 3612
rect 676 800 704 3606
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1124 2848 1176 2854
rect 1124 2790 1176 2796
rect 1136 800 1164 2790
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1320 649 1348 2382
rect 1412 1873 1440 2926
rect 1398 1864 1454 1873
rect 1398 1799 1454 1808
rect 1596 800 1624 3334
rect 1688 2854 1716 5646
rect 1964 3058 1992 6802
rect 2424 6730 2452 7346
rect 2884 7002 2912 7414
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2332 4146 2360 5170
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 2148 800 2176 3130
rect 2332 2514 2360 4082
rect 2424 2990 2452 6666
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 6322 2820 6598
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2516 4826 2544 5170
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2608 4622 2636 5510
rect 3160 4622 3188 7278
rect 3252 6254 3280 7890
rect 3804 7750 3832 8230
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 6390 3372 7346
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3528 6322 3556 6666
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 5778 3280 6190
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3398 2728 4014
rect 3068 3534 3096 4422
rect 3160 4146 3188 4558
rect 3252 4146 3280 5714
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3240 4140 3292 4146
rect 3528 4128 3556 6258
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3620 5370 3648 5510
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3620 4690 3648 5306
rect 3804 5166 3832 7686
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3896 5098 3924 9318
rect 3988 8090 4016 13126
rect 4632 12986 4660 14214
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12238 4660 12582
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11830 4384 12038
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4632 7478 4660 8230
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 5914 4016 6734
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5370 4108 6938
rect 4632 6798 4660 7414
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3700 4140 3752 4146
rect 3528 4100 3700 4128
rect 3240 4082 3292 4088
rect 3700 4082 3752 4088
rect 3160 3602 3188 4082
rect 3976 4072 4028 4078
rect 4172 4026 4200 4558
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4146 4384 4422
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 3976 4014 4028 4020
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2700 3058 2728 3334
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2608 800 2636 2858
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 2884 2281 2912 2790
rect 3056 2304 3108 2310
rect 2870 2272 2926 2281
rect 3056 2246 3108 2252
rect 2870 2207 2926 2216
rect 2780 1488 2832 1494
rect 2778 1456 2780 1465
rect 2832 1456 2834 1465
rect 2778 1391 2834 1400
rect 3068 800 3096 2246
rect 3424 1216 3476 1222
rect 3424 1158 3476 1164
rect 3436 1057 3464 1158
rect 3422 1048 3478 1057
rect 3422 983 3478 992
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3528 241 3556 2790
rect 3620 800 3648 3946
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3534 3924 3878
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3712 2922 3740 3402
rect 3988 3097 4016 4014
rect 4080 3998 4200 4026
rect 4080 3194 4108 3998
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3346 4660 5170
rect 4724 4060 4752 20810
rect 5000 18086 5028 22066
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 8242 5028 18022
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 16250 5396 16458
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 10130 5120 15846
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13938 5396 14214
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5460 10266 5488 22170
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6196 21010 6224 21966
rect 6288 21894 6316 33934
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6748 16114 6776 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 7564 32224 7616 32230
rect 7564 32166 7616 32172
rect 7576 21146 7604 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 7748 30320 7800 30326
rect 7748 30262 7800 30268
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7116 20602 7144 20810
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5828 14482 5856 15914
rect 6748 15638 6776 16050
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 7024 15570 7052 15846
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 13530 5764 14214
rect 6288 13870 6316 14418
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5644 13190 5672 13466
rect 5828 13410 5856 13670
rect 5736 13382 5856 13410
rect 5736 13326 5764 13382
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5552 11762 5580 13126
rect 6288 12866 6316 13806
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 6288 12838 6592 12866
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 12170 5672 12582
rect 5736 12434 5764 12786
rect 6288 12782 6316 12838
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12442 6500 12718
rect 6564 12714 6592 12838
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6460 12436 6512 12442
rect 5736 12406 5856 12434
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5828 11558 5856 12406
rect 6460 12378 6512 12384
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11762 6132 12174
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11150 5856 11494
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5000 8214 5120 8242
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 6662 4844 7278
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4724 4032 4844 4060
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4172 3318 4660 3346
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3974 3088 4030 3097
rect 3974 3023 4030 3032
rect 3700 2916 3752 2922
rect 4172 2904 4200 3318
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 3700 2858 3752 2864
rect 4080 2876 4200 2904
rect 4080 2689 4108 2876
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4066 2680 4122 2689
rect 4214 2683 4522 2692
rect 4066 2615 4122 2624
rect 4632 1578 4660 2994
rect 4724 2446 4752 3878
rect 4816 3738 4844 4032
rect 5092 3942 5120 8214
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4540 1550 4660 1578
rect 4540 800 4568 1550
rect 5092 800 5120 2926
rect 5184 1494 5212 4558
rect 5276 4010 5304 6122
rect 5368 4554 5396 10066
rect 5644 9110 5672 10134
rect 6104 10062 6132 11698
rect 6840 11626 6868 13466
rect 7116 12434 7144 19382
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17202 7420 17478
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7300 16590 7328 17138
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7300 16454 7328 16526
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16046 7328 16390
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7392 15978 7420 16730
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 12646 7420 14962
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7116 12406 7236 12434
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5736 8566 5764 9998
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6380 9722 6408 9930
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9178 5856 9318
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5920 8498 5948 8774
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5920 7546 5948 8434
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6012 7410 6040 9114
rect 6104 9110 6132 9522
rect 6196 9178 6224 9522
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6564 7886 6592 9930
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 6798 5488 7210
rect 6012 7002 6040 7346
rect 6564 7206 6592 7822
rect 6932 7410 6960 8502
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 7116 7546 7144 7754
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5460 5234 5488 6734
rect 6012 6390 6040 6734
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 6564 5778 6592 7142
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4758 5488 5170
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5736 3058 5764 4966
rect 6196 3126 6224 5510
rect 6564 4690 6592 5714
rect 6748 5574 6776 6802
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 5710 6868 6598
rect 7208 6254 7236 12406
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6798 7328 7346
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7392 6746 7420 12582
rect 7484 7478 7512 20538
rect 7576 19922 7604 21082
rect 7668 20448 7696 29174
rect 7760 21078 7788 30262
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 7748 21072 7800 21078
rect 7748 21014 7800 21020
rect 8036 20602 8064 21898
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8128 21010 8156 21830
rect 9692 21554 9720 21966
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10428 21146 10456 21490
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7668 20420 7788 20448
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7668 19378 7696 20266
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18766 7696 19314
rect 7760 18834 7788 20420
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 20058 7880 20334
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 8312 19854 8340 20878
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 20602 8432 20742
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8312 19378 8340 19790
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7668 18290 7696 18702
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7576 15026 7604 18158
rect 7668 17678 7696 18226
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17338 7696 17478
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15502 7696 16050
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12102 7696 12786
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11762 7696 12038
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7760 9738 7788 17682
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 16250 7880 16390
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 12434 7972 18702
rect 8312 18630 8340 19314
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8404 18902 8432 19246
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7852 12406 7972 12434
rect 7852 10146 7880 12406
rect 7852 10118 7972 10146
rect 7668 9710 7788 9738
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7668 6934 7696 9710
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7760 8566 7788 8978
rect 7852 8974 7880 9454
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7760 8090 7788 8502
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7410 7880 8910
rect 7944 7546 7972 10118
rect 8036 9586 8064 16050
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 12434 8248 15438
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15094 8340 15370
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8128 12406 8248 12434
rect 8128 10418 8156 12406
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8128 10390 8248 10418
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8128 8566 8156 9998
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8128 8294 8156 8502
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8220 7954 8248 10390
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 8022 8340 8230
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 7002 7880 7346
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7656 6792 7708 6798
rect 7392 6740 7656 6746
rect 7392 6734 7708 6740
rect 7392 6718 7696 6734
rect 7392 6390 7420 6718
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3534 6500 3878
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6288 3126 6316 3334
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6380 2990 6408 3334
rect 6564 3058 6592 4626
rect 6840 4146 6868 5238
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5644 2582 5672 2858
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 6380 2446 6408 2790
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 5172 1488 5224 1494
rect 5172 1430 5224 1436
rect 5552 800 5580 2382
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6012 800 6040 2246
rect 6472 800 6500 2450
rect 7116 1222 7144 3470
rect 7104 1216 7156 1222
rect 7104 1158 7156 1164
rect 7484 800 7512 3470
rect 7944 3194 7972 4150
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8220 3058 8248 4966
rect 8404 3942 8432 10950
rect 8496 10674 8524 14010
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8588 7818 8616 20402
rect 9416 19990 9444 21082
rect 10980 21078 11008 21286
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9416 19378 9444 19926
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18698 8708 19110
rect 9692 18766 9720 19246
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 9692 16590 9720 18702
rect 9784 18222 9812 19110
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9784 17202 9812 18158
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9232 14414 9260 14758
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8772 12850 8800 14350
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8772 12238 8800 12786
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 9324 11762 9352 16526
rect 9692 13326 9720 16526
rect 9784 13870 9812 17138
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9416 13190 9444 13262
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12986 9444 13126
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8680 11150 8708 11698
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9784 11150 9812 11562
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 8680 10674 8708 11086
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8680 10266 8708 10610
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9450 8892 9862
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8680 8498 8708 8910
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8680 7410 8708 8434
rect 8864 7410 8892 9386
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8864 6866 8892 7346
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 9324 3058 9352 11018
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 3738 9628 10406
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 5234 9812 7278
rect 9968 5914 9996 20946
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10152 18086 10180 18702
rect 10612 18426 10640 20878
rect 10980 20806 11008 20878
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 18766 11008 20742
rect 12268 19242 12296 25230
rect 13096 21146 13124 27406
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 15752 26444 15804 26450
rect 15752 26386 15804 26392
rect 15764 21146 15792 26386
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12544 20466 12572 20878
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19378 12388 19790
rect 12544 19446 12572 20402
rect 12728 20058 12756 20402
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12544 18766 12572 19382
rect 12820 19174 12848 19926
rect 13096 19854 13124 21082
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20602 14688 20810
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18970 12848 19110
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 12820 18290 12848 18906
rect 12912 18630 12940 19246
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13188 18766 13216 19110
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 16658 10180 18022
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10244 16522 10272 17138
rect 11520 17128 11572 17134
rect 11520 17070 11572 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10244 16114 10272 16458
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10336 15910 10364 16934
rect 11532 16794 11560 17070
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 12360 16590 12388 16934
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10980 15502 11008 16526
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15502 11192 15846
rect 11624 15638 11652 16050
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 10980 15094 11008 15438
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14618 10364 14826
rect 11256 14618 11284 14894
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 10520 13870 10548 14554
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 9586 10088 13262
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10152 12442 10180 12786
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 9580 10100 9586
rect 10048 9522 10100 9528
rect 10244 9042 10272 13806
rect 10520 13530 10548 13806
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10520 13394 10548 13466
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10888 13326 10916 14350
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 12238 10364 12582
rect 10520 12238 10548 13126
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 10336 11830 10364 12174
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 6798 10088 8842
rect 10244 8498 10272 8978
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 7886 10364 9454
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 8090 10548 8366
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10520 7206 10548 8026
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7410 10640 7686
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 10060 5166 10088 6734
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10520 6662 10548 7142
rect 10612 6662 10640 7346
rect 10796 7342 10824 7822
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10888 7290 10916 11018
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 7886 11008 9114
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 7954 11192 8570
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10888 7262 11008 7290
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9876 4826 9904 5102
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 10060 4622 10088 5102
rect 10520 5098 10548 6598
rect 10888 6458 10916 7142
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5370 10732 6122
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10704 5234 10732 5306
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4146 9812 4490
rect 10152 4282 10180 4966
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4282 10272 4422
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9048 2446 9076 2790
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 800 7972 2246
rect 8496 800 8524 2382
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 800 8984 2246
rect 9416 800 9444 2790
rect 10244 2650 10272 4082
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10428 800 10456 3470
rect 10796 3058 10824 3538
rect 10888 3194 10916 6258
rect 10980 4010 11008 7262
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4826 11192 5170
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 4146 11284 11494
rect 11716 11286 11744 12174
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 9450 11468 10542
rect 11992 10062 12020 11494
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12084 10266 12112 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11440 8974 11468 9386
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11440 8430 11468 8910
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8634 11560 8842
rect 11992 8634 12020 9998
rect 12176 8906 12204 15438
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 9110 12296 14962
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12728 13938 12756 14010
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12912 13326 12940 14350
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12442 12388 12854
rect 12912 12850 12940 13262
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 13188 12442 13216 13262
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 12716 12232 12768 12238
rect 12636 12180 12716 12186
rect 12636 12174 12768 12180
rect 12636 12158 12756 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11898 12572 12038
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 9926 12480 10950
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12544 9450 12572 11222
rect 12636 11150 12664 12158
rect 13188 11354 13216 12378
rect 13280 12374 13308 18702
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13464 18086 13492 18634
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13464 16182 13492 18022
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13464 16046 13492 16118
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13360 14340 13412 14346
rect 13360 14282 13412 14288
rect 13372 13326 13400 14282
rect 13464 14074 13492 15982
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13372 12238 13400 12718
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13372 11558 13400 11698
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12820 10810 12848 11086
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 13188 8566 13216 8774
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11716 6390 11744 8434
rect 11900 8090 11928 8434
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11348 4622 11376 6326
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4622 11560 4966
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11348 4078 11376 4558
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 11624 3738 11652 4558
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10980 3058 11008 3334
rect 11440 3058 11468 3470
rect 11900 3466 11928 3878
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11992 3194 12020 8434
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 8022 13124 8230
rect 13372 8090 13400 8910
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13084 8016 13136 8022
rect 13084 7958 13136 7964
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7342 13124 7686
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13188 7002 13216 7346
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13464 6390 13492 12310
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13556 5370 13584 20402
rect 15028 20058 15056 20402
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 19378 14688 19790
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18970 13768 19110
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 14292 18766 14320 19314
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17882 14412 18226
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14752 17610 14780 18566
rect 14936 18426 14964 18770
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13648 14278 13676 17002
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 15026 14228 15642
rect 14660 15638 14688 15846
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13924 13734 13952 14894
rect 14476 14414 14504 15438
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14292 13938 14320 14350
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13394 13952 13670
rect 14108 13530 14136 13874
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 12714 13768 13262
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11898 13676 12038
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 14660 11830 14688 12854
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7546 13860 7686
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7274 13860 7346
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 6322 13860 7210
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 10612 2446 10640 2994
rect 10796 2446 10824 2994
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10888 800 10916 2246
rect 11348 800 11376 2790
rect 11992 2446 12020 2858
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 800 11928 2246
rect 12360 800 12388 3470
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12636 3126 12664 3334
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12728 3058 12756 3334
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 13372 800 13400 3470
rect 14016 3194 14044 9998
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7206 14412 7686
rect 14476 7546 14504 8230
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14384 2650 14412 7142
rect 14476 6866 14504 7482
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14568 6458 14596 6734
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 2774 14688 7346
rect 14844 4826 14872 17614
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13258 15056 13670
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3058 14780 3470
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14568 2746 14688 2774
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13832 800 13860 2246
rect 14292 800 14320 2382
rect 14568 2106 14596 2746
rect 14844 2446 14872 3878
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3058 14964 3334
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14844 800 14872 2246
rect 15028 1970 15056 5646
rect 15120 5370 15148 20402
rect 15764 19854 15792 21082
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15212 5914 15240 19382
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18766 15608 19110
rect 16868 18970 16896 19246
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15304 17338 15332 18294
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15488 16726 15516 17478
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15488 16114 15516 16662
rect 16316 16658 16344 17274
rect 16684 17202 16712 17614
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15488 14482 15516 16050
rect 15672 15706 15700 16050
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12238 15332 12786
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 12442 15424 12582
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15304 11762 15332 12174
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15396 11558 15424 12378
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15580 8634 15608 13262
rect 15764 12434 15792 16050
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12986 15884 13126
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15856 12850 15884 12922
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15764 12406 15884 12434
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15672 10810 15700 11834
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 8634 15792 9522
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6866 15792 7142
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15304 5642 15332 6394
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15672 5710 15700 6326
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15304 5302 15332 5578
rect 15396 5574 15424 5646
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15396 5234 15424 5510
rect 15856 5370 15884 12406
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 11354 15976 11630
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16040 9178 16068 9522
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16132 8974 16160 9318
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15948 6798 15976 8434
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15016 1964 15068 1970
rect 15016 1906 15068 1912
rect 15120 1902 15148 5170
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15212 3058 15240 3402
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15304 800 15332 2450
rect 15672 2038 15700 5170
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15764 3126 15792 3606
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15660 2032 15712 2038
rect 15660 1974 15712 1980
rect 15856 1630 15884 4558
rect 15948 2378 15976 5646
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15844 1624 15896 1630
rect 15844 1566 15896 1572
rect 16040 1426 16068 6258
rect 16132 3670 16160 8434
rect 16224 8362 16252 16526
rect 16500 15910 16528 16730
rect 16960 16574 16988 17138
rect 17236 16794 17264 17546
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 16960 16546 17080 16574
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16684 16114 16712 16458
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16500 15638 16528 15846
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16500 14618 16528 15574
rect 16684 15502 16712 16050
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16684 14414 16712 15438
rect 17052 14958 17080 16546
rect 17328 15502 17356 21558
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 18064 17882 18092 19722
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 16250 17448 16390
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 14278 16896 14350
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 14074 16896 14214
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 12782 16896 13670
rect 16960 13530 16988 13874
rect 17052 13734 17080 14894
rect 17512 14618 17540 14962
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17236 13326 17264 14214
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12918 17172 13194
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16500 7954 16528 9454
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6390 16252 6734
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16316 4622 16344 6666
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16408 5914 16436 6258
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16500 5846 16528 7890
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 4078 16344 4558
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16316 3602 16344 4014
rect 16592 3738 16620 10610
rect 16684 8498 16712 12106
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16776 5658 16804 11766
rect 16868 11150 16896 12718
rect 16960 12442 16988 12786
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17144 12238 17172 12854
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12238 17356 12582
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 9382 16896 11086
rect 17144 10742 17172 12174
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 6186 16896 9318
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7342 17172 7822
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17144 6866 17172 7278
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16684 5630 16804 5658
rect 16684 4434 16712 5630
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5302 16804 5510
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16776 4554 16804 5238
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 16868 4690 16896 5170
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16684 4406 16804 4434
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16028 1420 16080 1426
rect 16028 1362 16080 1368
rect 16224 800 16252 3470
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 2854 16712 3334
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16776 2514 16804 4406
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16764 2508 16816 2514
rect 16764 2450 16816 2456
rect 16868 1442 16896 2790
rect 16960 2446 16988 3538
rect 17144 3398 17172 5170
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17052 2990 17080 3334
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17052 2774 17080 2926
rect 17052 2746 17172 2774
rect 17144 2446 17172 2746
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 16776 1414 16896 1442
rect 16776 800 16804 1414
rect 17236 800 17264 2246
rect 17328 1766 17356 8434
rect 17420 3194 17448 12174
rect 17512 3738 17540 13262
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 10810 17632 11018
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17788 5370 17816 16526
rect 18064 16114 18092 17818
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16794 18184 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 14414 17908 15302
rect 17972 15162 18000 15438
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17880 10810 17908 11494
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 7954 17908 8910
rect 18064 8838 18092 9318
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8566 18092 8774
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 18248 4826 18276 14350
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18432 6934 18460 7142
rect 18420 6928 18472 6934
rect 18420 6870 18472 6876
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 4214 18552 4422
rect 18512 4208 18564 4214
rect 18512 4150 18564 4156
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17604 3602 17632 4014
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17604 3058 17632 3538
rect 18524 3534 18552 4150
rect 18616 4146 18644 16526
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18708 11354 18736 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19260 9178 19288 9590
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19076 8634 19104 8842
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18800 7546 18828 8502
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5302 18920 6054
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18800 4690 18828 5170
rect 18892 4690 18920 5238
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18800 4146 18828 4626
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18340 3194 18368 3470
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 17684 2916 17736 2922
rect 17684 2858 17736 2864
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17604 1306 17632 2518
rect 17696 2446 17724 2858
rect 17972 2514 18000 2858
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17604 1278 17724 1306
rect 17696 800 17724 1278
rect 18708 800 18736 2926
rect 18984 2582 19012 2994
rect 19076 2650 19104 4558
rect 19168 3126 19196 8910
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19168 800 19196 2382
rect 19260 1494 19288 7346
rect 19352 5386 19380 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 19444 8498 19472 8910
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8566 20024 8774
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19444 7886 19472 8434
rect 19996 7954 20024 8502
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19352 5358 19472 5386
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19352 4554 19380 5238
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19444 4146 19472 5358
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19720 3602 19748 4082
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 2990 20024 3334
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19444 2446 19472 2790
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19248 1488 19300 1494
rect 19248 1430 19300 1436
rect 19720 870 19840 898
rect 19720 800 19748 870
rect 3514 232 3570 241
rect 3514 167 3570 176
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15750 0 15806 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 19812 762 19840 870
rect 19996 762 20024 2246
rect 20088 2038 20116 2246
rect 20076 2032 20128 2038
rect 20076 1974 20128 1980
rect 20180 800 20208 2790
rect 20456 1562 20484 8434
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20548 1698 20576 7822
rect 20640 1834 20668 8910
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20824 2038 20852 8434
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37280 6928 37332 6934
rect 37280 6870 37332 6876
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24596 4282 24624 4558
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24584 4276 24636 4282
rect 24584 4218 24636 4224
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21284 3058 21312 3946
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 21640 2848 21692 2854
rect 21640 2790 21692 2796
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 20812 2032 20864 2038
rect 20812 1974 20864 1980
rect 20628 1828 20680 1834
rect 20628 1770 20680 1776
rect 20536 1692 20588 1698
rect 20536 1634 20588 1640
rect 20444 1556 20496 1562
rect 20444 1498 20496 1504
rect 21100 800 21128 2382
rect 21192 2378 21220 2518
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21468 2106 21496 2450
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21560 2106 21588 2382
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 21548 2100 21600 2106
rect 21548 2042 21600 2048
rect 21652 800 21680 2790
rect 22204 2446 22232 2858
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 22112 800 22140 2246
rect 22572 800 22600 2382
rect 23584 800 23612 2994
rect 24688 2446 24716 4422
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24044 800 24072 2382
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24596 800 24624 2246
rect 25056 800 25084 2790
rect 25608 2650 25636 4082
rect 28816 4072 28868 4078
rect 28816 4014 28868 4020
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25700 2650 25728 3470
rect 28828 2650 28856 4014
rect 30300 2650 30328 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33324 2984 33376 2990
rect 33324 2926 33376 2932
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 25320 2576 25372 2582
rect 25320 2518 25372 2524
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 25332 2310 25360 2518
rect 25964 2440 26016 2446
rect 25964 2382 26016 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27988 2440 28040 2446
rect 27988 2382 28040 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 25976 800 26004 2382
rect 26528 800 26556 2382
rect 27448 800 27476 2382
rect 28000 800 28028 2382
rect 28920 800 28948 2382
rect 29472 800 29500 2382
rect 30392 800 30420 2382
rect 30484 1834 30512 2518
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31852 2440 31904 2446
rect 31852 2382 31904 2388
rect 30472 1828 30524 1834
rect 30472 1770 30524 1776
rect 30852 800 30880 2382
rect 31864 800 31892 2382
rect 32324 800 32352 2790
rect 33336 800 33364 2926
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 33796 800 33824 2382
rect 34808 800 34836 2382
rect 35176 1630 35204 2382
rect 35164 1624 35216 1630
rect 35164 1566 35216 1572
rect 35360 1442 35388 2790
rect 36268 2372 36320 2378
rect 36268 2314 36320 2320
rect 35268 1414 35388 1442
rect 35268 800 35296 1414
rect 36280 800 36308 2314
rect 36740 800 36768 2790
rect 37292 2650 37320 6870
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 38568 6316 38620 6322
rect 38568 6258 38620 6264
rect 37280 2644 37332 2650
rect 37280 2586 37332 2592
rect 38200 2440 38252 2446
rect 38200 2382 38252 2388
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37752 800 37780 2314
rect 38212 800 38240 2382
rect 38580 2378 38608 6258
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 59636 3460 59688 3466
rect 59636 3402 59688 3408
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 56692 3052 56744 3058
rect 56692 2994 56744 3000
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 42616 2848 42668 2854
rect 42616 2790 42668 2796
rect 44088 2848 44140 2854
rect 44088 2790 44140 2796
rect 46940 2848 46992 2854
rect 46940 2790 46992 2796
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 52828 2848 52880 2854
rect 52828 2790 52880 2796
rect 54300 2848 54352 2854
rect 54300 2790 54352 2796
rect 38568 2372 38620 2378
rect 38568 2314 38620 2320
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 39224 800 39252 2314
rect 39684 800 39712 2790
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 40408 2304 40460 2310
rect 40408 2246 40460 2252
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 40420 1902 40448 2246
rect 40408 1896 40460 1902
rect 40408 1838 40460 1844
rect 40512 1426 40540 2246
rect 40500 1420 40552 1426
rect 40500 1362 40552 1368
rect 40604 800 40632 2314
rect 41340 1306 41368 2382
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 41156 1278 41368 1306
rect 41156 800 41184 1278
rect 42076 800 42104 2314
rect 42628 800 42656 2790
rect 43076 2440 43128 2446
rect 43076 2382 43128 2388
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43088 1970 43116 2382
rect 43076 1964 43128 1970
rect 43076 1906 43128 1912
rect 43548 800 43576 2382
rect 44100 800 44128 2790
rect 45008 2440 45060 2446
rect 45008 2382 45060 2388
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 46480 2440 46532 2446
rect 46480 2382 46532 2388
rect 45020 800 45048 2382
rect 45480 800 45508 2382
rect 46492 800 46520 2382
rect 46756 2304 46808 2310
rect 46756 2246 46808 2252
rect 46768 2106 46796 2246
rect 46756 2100 46808 2106
rect 46756 2042 46808 2048
rect 46952 800 46980 2790
rect 47952 2440 48004 2446
rect 47952 2382 48004 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 49424 2440 49476 2446
rect 49424 2382 49476 2388
rect 47964 800 47992 2382
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 48332 1494 48360 2246
rect 48320 1488 48372 1494
rect 48320 1430 48372 1436
rect 48424 800 48452 2382
rect 49436 800 49464 2382
rect 49896 800 49924 2790
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 51356 2440 51408 2446
rect 51356 2382 51408 2388
rect 52368 2440 52420 2446
rect 52368 2382 52420 2388
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50908 800 50936 2382
rect 51172 2304 51224 2310
rect 51172 2246 51224 2252
rect 51184 2038 51212 2246
rect 51172 2032 51224 2038
rect 51172 1974 51224 1980
rect 51368 800 51396 2382
rect 52380 800 52408 2382
rect 52840 800 52868 2790
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 52920 2304 52972 2310
rect 52920 2246 52972 2252
rect 52932 1562 52960 2246
rect 52920 1556 52972 1562
rect 52920 1498 52972 1504
rect 53852 800 53880 2382
rect 54312 800 54340 2790
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 55772 2440 55824 2446
rect 55772 2382 55824 2388
rect 55232 800 55260 2382
rect 55496 2304 55548 2310
rect 55496 2246 55548 2252
rect 55508 1698 55536 2246
rect 55496 1692 55548 1698
rect 55496 1634 55548 1640
rect 55784 800 55812 2382
rect 56704 800 56732 2994
rect 58716 2848 58768 2854
rect 58716 2790 58768 2796
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 57060 2304 57112 2310
rect 57060 2246 57112 2252
rect 57072 1766 57100 2246
rect 57060 1760 57112 1766
rect 57060 1702 57112 1708
rect 57256 800 57284 2382
rect 58164 2372 58216 2378
rect 58164 2314 58216 2320
rect 58176 800 58204 2314
rect 58728 800 58756 2790
rect 59648 800 59676 3402
rect 19812 734 20024 762
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24030 0 24086 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39210 0 39266 800
rect 39670 0 39726 800
rect 40130 0 40186 800
rect 40590 0 40646 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50894 0 50950 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
<< via2 >>
rect 2778 41656 2834 41712
rect 1582 40840 1638 40896
rect 1490 40024 1546 40080
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 1582 38392 1638 38448
rect 1398 26560 1454 26616
rect 1582 37612 1584 37632
rect 1584 37612 1636 37632
rect 1636 37612 1638 37632
rect 1582 37576 1638 37612
rect 1582 36644 1638 36680
rect 1582 36624 1584 36644
rect 1584 36624 1636 36644
rect 1636 36624 1638 36644
rect 1582 35808 1638 35864
rect 1582 34992 1638 35048
rect 1582 34176 1638 34232
rect 1582 33804 1584 33824
rect 1584 33804 1636 33824
rect 1636 33804 1638 33824
rect 1582 33768 1638 33804
rect 1582 32952 1638 33008
rect 1582 32408 1638 32464
rect 1582 31592 1638 31648
rect 1582 31204 1638 31240
rect 1582 31184 1584 31204
rect 1584 31184 1636 31204
rect 1636 31184 1638 31204
rect 1582 30368 1638 30424
rect 1582 29996 1584 30016
rect 1584 29996 1636 30016
rect 1636 29996 1638 30016
rect 1582 29960 1638 29996
rect 1582 29144 1638 29200
rect 1582 28736 1638 28792
rect 1582 27376 1638 27432
rect 1582 26188 1584 26208
rect 1584 26188 1636 26208
rect 1636 26188 1638 26208
rect 1582 26152 1638 26188
rect 1582 25336 1638 25392
rect 1582 24928 1638 24984
rect 1582 24112 1638 24168
rect 1582 23704 1638 23760
rect 1582 22752 1638 22808
rect 1398 21528 1454 21584
rect 1398 20304 1454 20360
rect 1398 16496 1454 16552
rect 1582 22380 1584 22400
rect 1584 22380 1636 22400
rect 1636 22380 1638 22400
rect 1582 22344 1638 22380
rect 1582 21120 1638 21176
rect 1582 19932 1584 19952
rect 1584 19932 1636 19952
rect 1636 19932 1638 19952
rect 1582 19896 1638 19932
rect 1582 18572 1584 18592
rect 1584 18572 1636 18592
rect 1636 18572 1638 18592
rect 1582 18536 1638 18572
rect 1582 17720 1638 17776
rect 1582 17332 1638 17368
rect 1582 17312 1584 17332
rect 1584 17312 1636 17332
rect 1636 17312 1638 17332
rect 1582 16088 1638 16144
rect 1582 15272 1638 15328
rect 1582 14884 1638 14920
rect 1582 14864 1584 14884
rect 1584 14864 1636 14884
rect 1636 14864 1638 14884
rect 1582 13912 1638 13968
rect 1582 13524 1638 13560
rect 1582 13504 1584 13524
rect 1584 13504 1636 13524
rect 1636 13504 1638 13524
rect 1398 12688 1454 12744
rect 1582 12280 1638 12336
rect 3054 39244 3056 39264
rect 3056 39244 3108 39264
rect 3108 39244 3110 39264
rect 3054 39208 3110 39244
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2226 19080 2282 19136
rect 3054 27784 3110 27840
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1398 11464 1454 11520
rect 1582 11056 1638 11112
rect 1398 9832 1454 9888
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 2778 10240 2834 10296
rect 1582 8472 1638 8528
rect 2778 8064 2834 8120
rect 1582 7692 1584 7712
rect 1584 7692 1636 7712
rect 1636 7692 1638 7712
rect 1582 7656 1638 7692
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1490 6840 1546 6896
rect 1398 6432 1454 6488
rect 1582 6060 1584 6080
rect 1584 6060 1636 6080
rect 1636 6060 1638 6080
rect 1582 6024 1638 6060
rect 1582 4664 1638 4720
rect 1582 4256 1638 4312
rect 1398 1808 1454 1864
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 2870 2216 2926 2272
rect 2778 1436 2780 1456
rect 2780 1436 2832 1456
rect 2832 1436 2834 1456
rect 2778 1400 2834 1436
rect 3422 992 3478 1048
rect 1306 584 1362 640
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 3974 3032 4030 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2624 4122 2680
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 3514 176 3570 232
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 0 41714 800 41744
rect 2773 41714 2839 41717
rect 0 41712 2839 41714
rect 0 41656 2778 41712
rect 2834 41656 2839 41712
rect 0 41654 2839 41656
rect 0 41624 800 41654
rect 2773 41651 2839 41654
rect 0 41216 800 41336
rect 0 40898 800 40928
rect 1577 40898 1643 40901
rect 0 40896 1643 40898
rect 0 40840 1582 40896
rect 1638 40840 1643 40896
rect 0 40838 1643 40840
rect 0 40808 800 40838
rect 1577 40835 1643 40838
rect 0 40400 800 40520
rect 0 40082 800 40112
rect 1485 40082 1551 40085
rect 0 40080 1551 40082
rect 0 40024 1490 40080
rect 1546 40024 1551 40080
rect 0 40022 1551 40024
rect 0 39992 800 40022
rect 1485 40019 1551 40022
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39266 800 39296
rect 3049 39266 3115 39269
rect 0 39264 3115 39266
rect 0 39208 3054 39264
rect 3110 39208 3115 39264
rect 0 39206 3115 39208
rect 0 39176 800 39206
rect 3049 39203 3115 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 0 38768 800 38888
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38450 800 38480
rect 1577 38450 1643 38453
rect 0 38448 1643 38450
rect 0 38392 1582 38448
rect 1638 38392 1643 38448
rect 0 38390 1643 38392
rect 0 38360 800 38390
rect 1577 38387 1643 38390
rect 19570 38112 19886 38113
rect 0 37952 800 38072
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37634 800 37664
rect 1577 37634 1643 37637
rect 0 37632 1643 37634
rect 0 37576 1582 37632
rect 1638 37576 1643 37632
rect 0 37574 1643 37576
rect 0 37544 800 37574
rect 1577 37571 1643 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 0 37000 800 37120
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36682 800 36712
rect 1577 36682 1643 36685
rect 0 36680 1643 36682
rect 0 36624 1582 36680
rect 1638 36624 1643 36680
rect 0 36622 1643 36624
rect 0 36592 800 36622
rect 1577 36619 1643 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36184 800 36304
rect 19570 35936 19886 35937
rect 0 35866 800 35896
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 1577 35866 1643 35869
rect 0 35864 1643 35866
rect 0 35808 1582 35864
rect 1638 35808 1643 35864
rect 0 35806 1643 35808
rect 0 35776 800 35806
rect 1577 35803 1643 35806
rect 0 35368 800 35488
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 0 34552 800 34672
rect 4210 34304 4526 34305
rect 0 34234 800 34264
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 1577 34234 1643 34237
rect 0 34232 1643 34234
rect 0 34176 1582 34232
rect 1638 34176 1643 34232
rect 0 34174 1643 34176
rect 0 34144 800 34174
rect 1577 34171 1643 34174
rect 0 33826 800 33856
rect 1577 33826 1643 33829
rect 0 33824 1643 33826
rect 0 33768 1582 33824
rect 1638 33768 1643 33824
rect 0 33766 1643 33768
rect 0 33736 800 33766
rect 1577 33763 1643 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 0 33328 800 33448
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 33010 800 33040
rect 1577 33010 1643 33013
rect 0 33008 1643 33010
rect 0 32952 1582 33008
rect 1638 32952 1643 33008
rect 0 32950 1643 32952
rect 0 32920 800 32950
rect 1577 32947 1643 32950
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4210 32128 4526 32129
rect 0 31968 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 0 31650 800 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 800 31590
rect 1577 31587 1643 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 1577 31242 1643 31245
rect 0 31240 1643 31242
rect 0 31184 1582 31240
rect 1638 31184 1643 31240
rect 0 31182 1643 31184
rect 0 31152 800 31182
rect 1577 31179 1643 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30744 800 30864
rect 19570 30496 19886 30497
rect 0 30426 800 30456
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 1577 30426 1643 30429
rect 0 30424 1643 30426
rect 0 30368 1582 30424
rect 1638 30368 1643 30424
rect 0 30366 1643 30368
rect 0 30336 800 30366
rect 1577 30363 1643 30366
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 0 29520 800 29640
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 0 29202 800 29232
rect 1577 29202 1643 29205
rect 0 29200 1643 29202
rect 0 29144 1582 29200
rect 1638 29144 1643 29200
rect 0 29142 1643 29144
rect 0 29112 800 29142
rect 1577 29139 1643 29142
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 1577 28794 1643 28797
rect 0 28792 1643 28794
rect 0 28736 1582 28792
rect 1638 28736 1643 28792
rect 0 28734 1643 28736
rect 0 28704 800 28734
rect 1577 28731 1643 28734
rect 0 28296 800 28416
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 27842 800 27872
rect 3049 27842 3115 27845
rect 0 27840 3115 27842
rect 0 27784 3054 27840
rect 3110 27784 3115 27840
rect 0 27782 3115 27784
rect 0 27752 800 27782
rect 3049 27779 3115 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27434 800 27464
rect 1577 27434 1643 27437
rect 0 27432 1643 27434
rect 0 27376 1582 27432
rect 1638 27376 1643 27432
rect 0 27374 1643 27376
rect 0 27344 800 27374
rect 1577 27371 1643 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 0 26936 800 27056
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1393 26618 1459 26621
rect 0 26616 1459 26618
rect 0 26560 1398 26616
rect 1454 26560 1459 26616
rect 0 26558 1459 26560
rect 0 26528 800 26558
rect 1393 26555 1459 26558
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 0 25712 800 25832
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25394 800 25424
rect 1577 25394 1643 25397
rect 0 25392 1643 25394
rect 0 25336 1582 25392
rect 1638 25336 1643 25392
rect 0 25334 1643 25336
rect 0 25304 800 25334
rect 1577 25331 1643 25334
rect 19570 25056 19886 25057
rect 0 24986 800 25016
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 800 24926
rect 1577 24923 1643 24926
rect 0 24488 800 24608
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 0 23762 800 23792
rect 1577 23762 1643 23765
rect 0 23760 1643 23762
rect 0 23704 1582 23760
rect 1638 23704 1643 23760
rect 0 23702 1643 23704
rect 0 23672 800 23702
rect 1577 23699 1643 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23128 800 23248
rect 19570 22880 19886 22881
rect 0 22810 800 22840
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 1577 22810 1643 22813
rect 0 22808 1643 22810
rect 0 22752 1582 22808
rect 1638 22752 1643 22808
rect 0 22750 1643 22752
rect 0 22720 800 22750
rect 1577 22747 1643 22750
rect 0 22402 800 22432
rect 1577 22402 1643 22405
rect 0 22400 1643 22402
rect 0 22344 1582 22400
rect 1638 22344 1643 22400
rect 0 22342 1643 22344
rect 0 22312 800 22342
rect 1577 22339 1643 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21904 800 22024
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21586 800 21616
rect 1393 21586 1459 21589
rect 0 21584 1459 21586
rect 0 21528 1398 21584
rect 1454 21528 1459 21584
rect 0 21526 1459 21528
rect 0 21496 800 21526
rect 1393 21523 1459 21526
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1577 21178 1643 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 0 20680 800 20800
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 0 20362 800 20392
rect 1393 20362 1459 20365
rect 0 20360 1459 20362
rect 0 20304 1398 20360
rect 1454 20304 1459 20360
rect 0 20302 1459 20304
rect 0 20272 800 20302
rect 1393 20299 1459 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19954 800 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 800 19894
rect 1577 19891 1643 19894
rect 19570 19616 19886 19617
rect 0 19456 800 19576
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 0 19138 800 19168
rect 2221 19138 2287 19141
rect 0 19136 2287 19138
rect 0 19080 2226 19136
rect 2282 19080 2287 19136
rect 0 19078 2287 19080
rect 0 19048 800 19078
rect 2221 19075 2287 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 0 18594 800 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 800 18534
rect 1577 18531 1643 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 0 18096 800 18216
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 800 17718
rect 1577 17715 1643 17718
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 0 16872 800 16992
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16554 800 16584
rect 1393 16554 1459 16557
rect 0 16552 1459 16554
rect 0 16496 1398 16552
rect 1454 16496 1459 16552
rect 0 16494 1459 16496
rect 0 16464 800 16494
rect 1393 16491 1459 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 0 14922 800 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 800 14862
rect 1577 14859 1643 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14424 800 14544
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 0 13970 800 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 800 13910
rect 1577 13907 1643 13910
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 1577 13562 1643 13565
rect 0 13560 1643 13562
rect 0 13504 1582 13560
rect 1638 13504 1643 13560
rect 0 13502 1643 13504
rect 0 13472 800 13502
rect 1577 13499 1643 13502
rect 0 13064 800 13184
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 0 12746 800 12776
rect 1393 12746 1459 12749
rect 0 12744 1459 12746
rect 0 12688 1398 12744
rect 1454 12688 1459 12744
rect 0 12686 1459 12688
rect 0 12656 800 12686
rect 1393 12683 1459 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 19570 12000 19886 12001
rect 0 11840 800 11960
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11522 800 11552
rect 1393 11522 1459 11525
rect 0 11520 1459 11522
rect 0 11464 1398 11520
rect 1454 11464 1459 11520
rect 0 11462 1459 11464
rect 0 11432 800 11462
rect 1393 11459 1459 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 11114 800 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 800 11054
rect 1577 11051 1643 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 0 10616 800 10736
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 0 9890 800 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 800 9830
rect 1393 9827 1459 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8848 800 8968
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8530 800 8560
rect 1577 8530 1643 8533
rect 0 8528 1643 8530
rect 0 8472 1582 8528
rect 1638 8472 1643 8528
rect 0 8470 1643 8472
rect 0 8440 800 8470
rect 1577 8467 1643 8470
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 800 8062
rect 2773 8059 2839 8062
rect 0 7714 800 7744
rect 1577 7714 1643 7717
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 0 7624 800 7654
rect 1577 7651 1643 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 0 7216 800 7336
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 19570 6560 19886 6561
rect 0 6490 800 6520
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 1393 6490 1459 6493
rect 0 6488 1459 6490
rect 0 6432 1398 6488
rect 1454 6432 1459 6488
rect 0 6430 1459 6432
rect 0 6400 800 6430
rect 1393 6427 1459 6430
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5584 800 5704
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5176 800 5296
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 0 4722 800 4752
rect 1577 4722 1643 4725
rect 0 4720 1643 4722
rect 0 4664 1582 4720
rect 1638 4664 1643 4720
rect 0 4662 1643 4664
rect 0 4632 800 4662
rect 1577 4659 1643 4662
rect 19570 4384 19886 4385
rect 0 4314 800 4344
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 1577 4314 1643 4317
rect 0 4312 1643 4314
rect 0 4256 1582 4312
rect 1638 4256 1643 4312
rect 0 4254 1643 4256
rect 0 4224 800 4254
rect 1577 4251 1643 4254
rect 0 3816 800 3936
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3408 800 3528
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 0 3090 800 3120
rect 3969 3090 4035 3093
rect 0 3088 4035 3090
rect 0 3032 3974 3088
rect 4030 3032 4035 3088
rect 0 3030 4035 3032
rect 0 3000 800 3030
rect 3969 3027 4035 3030
rect 4210 2752 4526 2753
rect 0 2682 800 2712
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4061 2682 4127 2685
rect 0 2680 4127 2682
rect 0 2624 4066 2680
rect 4122 2624 4127 2680
rect 0 2622 4127 2624
rect 0 2592 800 2622
rect 4061 2619 4127 2622
rect 0 2274 800 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 800 2214
rect 2865 2211 2931 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 0 1866 800 1896
rect 1393 1866 1459 1869
rect 0 1864 1459 1866
rect 0 1808 1398 1864
rect 1454 1808 1459 1864
rect 0 1806 1459 1808
rect 0 1776 800 1806
rect 1393 1803 1459 1806
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 0 1050 800 1080
rect 3417 1050 3483 1053
rect 0 1048 3483 1050
rect 0 992 3422 1048
rect 3478 992 3483 1048
rect 0 990 3483 992
rect 0 960 800 990
rect 3417 987 3483 990
rect 0 642 800 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 800 582
rect 1301 579 1367 582
rect 0 234 800 264
rect 3509 234 3575 237
rect 0 232 3575 234
rect 0 176 3514 232
rect 3570 176 3575 232
rect 0 174 3575 176
rect 0 144 800 174
rect 3509 171 3575 174
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 39200 19888 39760
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 39744 35248 39760
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 39200 50608 39760
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_19 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1644511149
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1644511149
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1644511149
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_160
timestamp 1644511149
transform 1 0 15824 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1644511149
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1644511149
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1644511149
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1644511149
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_244
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_260
timestamp 1644511149
transform 1 0 25024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1644511149
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_300
timestamp 1644511149
transform 1 0 28704 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_312
timestamp 1644511149
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_316
timestamp 1644511149
transform 1 0 30176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_347
timestamp 1644511149
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_355
timestamp 1644511149
transform 1 0 33764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1644511149
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1644511149
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1644511149
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1644511149
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1644511149
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1644511149
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1644511149
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1644511149
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1644511149
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_493
timestamp 1644511149
transform 1 0 46460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_509
timestamp 1644511149
transform 1 0 47932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_514
timestamp 1644511149
transform 1 0 48392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_521
timestamp 1644511149
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_537
timestamp 1644511149
transform 1 0 50508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_541
timestamp 1644511149
transform 1 0 50876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_546
timestamp 1644511149
transform 1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1644511149
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1644511149
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_565
timestamp 1644511149
transform 1 0 53084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1644511149
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1644511149
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1644511149
transform 1 0 55660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_600
timestamp 1644511149
transform 1 0 56304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1644511149
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1644511149
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_33
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1644511149
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1644511149
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_116
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_120
timestamp 1644511149
transform 1 0 12144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1644511149
transform 1 0 12788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1644511149
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_151
timestamp 1644511149
transform 1 0 14996 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1644511149
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1644511149
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_203
timestamp 1644511149
transform 1 0 19780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_207
timestamp 1644511149
transform 1 0 20148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_211
timestamp 1644511149
transform 1 0 20516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_228 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_260
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_264
timestamp 1644511149
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_343
timestamp 1644511149
transform 1 0 32660 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_369
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_375
timestamp 1644511149
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1644511149
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_396
timestamp 1644511149
transform 1 0 37536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_408
timestamp 1644511149
transform 1 0 38640 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_423
timestamp 1644511149
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_455
timestamp 1644511149
transform 1 0 42964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_467
timestamp 1644511149
transform 1 0 44068 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_471
timestamp 1644511149
transform 1 0 44436 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_483
timestamp 1644511149
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_508
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_520
timestamp 1644511149
transform 1 0 48944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_528
timestamp 1644511149
transform 1 0 49680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_534
timestamp 1644511149
transform 1 0 50232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_546
timestamp 1644511149
transform 1 0 51336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1644511149
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_566
timestamp 1644511149
transform 1 0 53176 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_578
timestamp 1644511149
transform 1 0 54280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_582
timestamp 1644511149
transform 1 0 54648 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_594
timestamp 1644511149
transform 1 0 55752 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_602
timestamp 1644511149
transform 1 0 56488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1644511149
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1644511149
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1644511149
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1644511149
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1644511149
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_116
timestamp 1644511149
transform 1 0 11776 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_126
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1644511149
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_174
timestamp 1644511149
transform 1 0 17112 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1644511149
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1644511149
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50
timestamp 1644511149
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_66
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_78
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1644511149
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_179
timestamp 1644511149
transform 1 0 17572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1644511149
transform 1 0 2300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1644511149
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_48
timestamp 1644511149
transform 1 0 5520 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_59
timestamp 1644511149
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_71
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_101
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1644511149
transform 1 0 11684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1644511149
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_207
timestamp 1644511149
transform 1 0 20148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_219
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_231
timestamp 1644511149
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1644511149
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_256
timestamp 1644511149
transform 1 0 24656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_268
timestamp 1644511149
transform 1 0 25760 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1644511149
transform 1 0 26864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_292
timestamp 1644511149
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_6
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1644511149
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1644511149
transform 1 0 6808 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1644511149
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_86
timestamp 1644511149
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1644511149
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1644511149
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1644511149
transform 1 0 12972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1644511149
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1644511149
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_175
timestamp 1644511149
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp 1644511149
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1644511149
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1644511149
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1644511149
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_56
timestamp 1644511149
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_151
timestamp 1644511149
transform 1 0 14996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_155
timestamp 1644511149
transform 1 0 15364 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_162
timestamp 1644511149
transform 1 0 16008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_187
timestamp 1644511149
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1644511149
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1644511149
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1644511149
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_92
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_100
timestamp 1644511149
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_107
timestamp 1644511149
transform 1 0 10948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_147
timestamp 1644511149
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1644511149
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_194
timestamp 1644511149
transform 1 0 18952 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_206
timestamp 1644511149
transform 1 0 20056 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1644511149
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1644511149
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1644511149
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_47
timestamp 1644511149
transform 1 0 5428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_71
timestamp 1644511149
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1644511149
transform 1 0 9568 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_96
timestamp 1644511149
transform 1 0 9936 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_113
timestamp 1644511149
transform 1 0 11500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_125
timestamp 1644511149
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1644511149
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_159
timestamp 1644511149
transform 1 0 15732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1644511149
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1644511149
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1644511149
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1644511149
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1644511149
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1644511149
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1644511149
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1644511149
transform 1 0 13248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1644511149
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1644511149
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_152
timestamp 1644511149
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_173
timestamp 1644511149
transform 1 0 17020 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1644511149
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_194
timestamp 1644511149
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_206
timestamp 1644511149
transform 1 0 20056 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1644511149
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_126
timestamp 1644511149
transform 1 0 12696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_203
timestamp 1644511149
transform 1 0 19780 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1644511149
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_10
timestamp 1644511149
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1644511149
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_60
timestamp 1644511149
transform 1 0 6624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_77
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_119
timestamp 1644511149
transform 1 0 12052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_127
timestamp 1644511149
transform 1 0 12788 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1644511149
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1644511149
transform 1 0 17204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1644511149
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_195
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1644511149
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_13
timestamp 1644511149
transform 1 0 2300 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp 1644511149
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1644511149
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_119
timestamp 1644511149
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1644511149
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1644511149
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_203
timestamp 1644511149
transform 1 0 19780 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1644511149
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1644511149
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1644511149
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_60
timestamp 1644511149
transform 1 0 6624 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_72
timestamp 1644511149
transform 1 0 7728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1644511149
transform 1 0 9016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1644511149
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_185
timestamp 1644511149
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_197
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_209
timestamp 1644511149
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1644511149
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1644511149
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1644511149
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_48
timestamp 1644511149
transform 1 0 5520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1644511149
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_125
timestamp 1644511149
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_25
timestamp 1644511149
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_77
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_85
timestamp 1644511149
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_97
timestamp 1644511149
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1644511149
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1644511149
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_153
timestamp 1644511149
transform 1 0 15180 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1644511149
transform 1 0 18032 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1644511149
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1644511149
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_14
timestamp 1644511149
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1644511149
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_162
timestamp 1644511149
transform 1 0 16008 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1644511149
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_24
timestamp 1644511149
transform 1 0 3312 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_83
timestamp 1644511149
transform 1 0 8740 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_95
timestamp 1644511149
transform 1 0 9844 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1644511149
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_121
timestamp 1644511149
transform 1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_129
timestamp 1644511149
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_138
timestamp 1644511149
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1644511149
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1644511149
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_201
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_213
timestamp 1644511149
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1644511149
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_6
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1644511149
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_38
timestamp 1644511149
transform 1 0 4600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_50
timestamp 1644511149
transform 1 0 5704 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_72
timestamp 1644511149
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1644511149
transform 1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_112
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1644511149
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1644511149
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_42
timestamp 1644511149
transform 1 0 4968 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_48
timestamp 1644511149
transform 1 0 5520 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1644511149
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1644511149
transform 1 0 7176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_78
timestamp 1644511149
transform 1 0 8280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1644511149
transform 1 0 8648 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1644511149
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_156
timestamp 1644511149
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_213
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1644511149
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1644511149
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1644511149
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_33
timestamp 1644511149
transform 1 0 4140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1644511149
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_63
timestamp 1644511149
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1644511149
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1644511149
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_108
timestamp 1644511149
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_120
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1644511149
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1644511149
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_33
timestamp 1644511149
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_45
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_152
timestamp 1644511149
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1644511149
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_6
timestamp 1644511149
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_12
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1644511149
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_37
timestamp 1644511149
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_45
timestamp 1644511149
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_55
timestamp 1644511149
transform 1 0 6164 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_67
timestamp 1644511149
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1644511149
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1644511149
transform 1 0 11316 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1644511149
transform 1 0 13156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_151
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_163
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1644511149
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1644511149
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1644511149
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_191
timestamp 1644511149
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1644511149
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_10
timestamp 1644511149
transform 1 0 2024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1644511149
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_62
timestamp 1644511149
transform 1 0 6808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1644511149
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1644511149
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_150
timestamp 1644511149
transform 1 0 14904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_162
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_174
timestamp 1644511149
transform 1 0 17112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1644511149
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_26
timestamp 1644511149
transform 1 0 3496 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_38
timestamp 1644511149
transform 1 0 4600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1644511149
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_75
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1644511149
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_130
timestamp 1644511149
transform 1 0 13064 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_150
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_178
timestamp 1644511149
transform 1 0 17480 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_202
timestamp 1644511149
transform 1 0 19688 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_214
timestamp 1644511149
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_49
timestamp 1644511149
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_61
timestamp 1644511149
transform 1 0 6716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_72
timestamp 1644511149
transform 1 0 7728 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1644511149
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_115
timestamp 1644511149
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1644511149
transform 1 0 12604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1644511149
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1644511149
transform 1 0 16836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1644511149
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_19
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_31
timestamp 1644511149
transform 1 0 3956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_43
timestamp 1644511149
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_72
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_84
timestamp 1644511149
transform 1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1644511149
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp 1644511149
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_211
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_49
timestamp 1644511149
transform 1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1644511149
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1644511149
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_150
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_162
timestamp 1644511149
transform 1 0 16008 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_168
timestamp 1644511149
transform 1 0 16560 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1644511149
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1644511149
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1644511149
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1644511149
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1644511149
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1644511149
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_7
timestamp 1644511149
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_48
timestamp 1644511149
transform 1 0 5520 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_60
timestamp 1644511149
transform 1 0 6624 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1644511149
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1644511149
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_89
timestamp 1644511149
transform 1 0 9292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_101
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1644511149
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_148
timestamp 1644511149
transform 1 0 14720 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_184
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_6
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_25
timestamp 1644511149
transform 1 0 3404 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1644511149
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1644511149
transform 1 0 6992 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_74
timestamp 1644511149
transform 1 0 7912 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_83
timestamp 1644511149
transform 1 0 8740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_97
timestamp 1644511149
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1644511149
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_132
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_144
timestamp 1644511149
transform 1 0 14352 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1644511149
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_74
timestamp 1644511149
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1644511149
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_164
timestamp 1644511149
transform 1 0 16192 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_176
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1644511149
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_25
timestamp 1644511149
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_37
timestamp 1644511149
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1644511149
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_121
timestamp 1644511149
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1644511149
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_6
timestamp 1644511149
transform 1 0 1656 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_33
timestamp 1644511149
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_44
timestamp 1644511149
transform 1 0 5152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_52
timestamp 1644511149
transform 1 0 5888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_71
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_95
timestamp 1644511149
transform 1 0 9844 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_107
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1644511149
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_160
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1644511149
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_25
timestamp 1644511149
transform 1 0 3404 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1644511149
transform 1 0 4048 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1644511149
transform 1 0 5152 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_89
timestamp 1644511149
transform 1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_33
timestamp 1644511149
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_40
timestamp 1644511149
transform 1 0 4784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_52
timestamp 1644511149
transform 1 0 5888 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1644511149
transform 1 0 3220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1644511149
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_41
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_6
timestamp 1644511149
transform 1 0 1656 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 1644511149
transform 1 0 2760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1644511149
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1644511149
transform 1 0 3036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1644511149
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1644511149
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_6
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_34
timestamp 1644511149
transform 1 0 4232 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_46
timestamp 1644511149
transform 1 0 5336 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1644511149
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1644511149
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_45
timestamp 1644511149
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_57
timestamp 1644511149
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1644511149
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_18
timestamp 1644511149
transform 1 0 2760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_26
timestamp 1644511149
transform 1 0 3496 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1644511149
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1644511149
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_21
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_35
timestamp 1644511149
transform 1 0 4324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_47
timestamp 1644511149
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_59
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_23
timestamp 1644511149
transform 1 0 3220 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_34
timestamp 1644511149
transform 1 0 4232 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1644511149
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1644511149
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_11
timestamp 1644511149
transform 1 0 2116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_49
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_6
timestamp 1644511149
transform 1 0 1656 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_12
timestamp 1644511149
transform 1 0 2208 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_16
timestamp 1644511149
transform 1 0 2576 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_24
timestamp 1644511149
transform 1 0 3312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_35
timestamp 1644511149
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1644511149
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_13
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_6
timestamp 1644511149
transform 1 0 1656 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_18
timestamp 1644511149
transform 1 0 2760 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1644511149
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_38
timestamp 1644511149
transform 1 0 4600 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_50
timestamp 1644511149
transform 1 0 5704 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_62
timestamp 1644511149
transform 1 0 6808 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_74
timestamp 1644511149
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1644511149
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_38
timestamp 1644511149
transform 1 0 4600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_50
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_6
timestamp 1644511149
transform 1 0 1656 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_14
timestamp 1644511149
transform 1 0 2392 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1644511149
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_35
timestamp 1644511149
transform 1 0 4324 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1644511149
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1644511149
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_22
timestamp 1644511149
transform 1 0 3128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_37
timestamp 1644511149
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_43
timestamp 1644511149
transform 1 0 5060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_55
timestamp 1644511149
transform 1 0 6164 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_67
timestamp 1644511149
transform 1 0 7268 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1644511149
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_7
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_13
timestamp 1644511149
transform 1 0 2300 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_23
timestamp 1644511149
transform 1 0 3220 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_35
timestamp 1644511149
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_46
timestamp 1644511149
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_58
timestamp 1644511149
transform 1 0 6440 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_70
timestamp 1644511149
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1644511149
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_6
timestamp 1644511149
transform 1 0 1656 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 1644511149
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1644511149
transform 1 0 1656 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1644511149
transform 1 0 2760 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1644511149
transform 1 0 3864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1644511149
transform 1 0 4968 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1644511149
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 1644511149
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_31
timestamp 1644511149
transform 1 0 3956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_43
timestamp 1644511149
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_513
timestamp 1644511149
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_569
timestamp 1644511149
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_7
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_31
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_43
timestamp 1644511149
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1644511149
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_517
timestamp 1644511149
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_529
timestamp 1644511149
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_541
timestamp 1644511149
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1644511149
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1644511149
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_561
timestamp 1644511149
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_573
timestamp 1644511149
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_585
timestamp 1644511149
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_597
timestamp 1644511149
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1644511149
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1644511149
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1644511149
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1644511149
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_513
timestamp 1644511149
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1644511149
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1644511149
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_533
timestamp 1644511149
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_545
timestamp 1644511149
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_557
timestamp 1644511149
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_569
timestamp 1644511149
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1644511149
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1644511149
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_589
timestamp 1644511149
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_601
timestamp 1644511149
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_613
timestamp 1644511149
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_7
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_19
timestamp 1644511149
transform 1 0 2852 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1644511149
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_517
timestamp 1644511149
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_529
timestamp 1644511149
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_541
timestamp 1644511149
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1644511149
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1644511149
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_561
timestamp 1644511149
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_573
timestamp 1644511149
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_585
timestamp 1644511149
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_597
timestamp 1644511149
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1644511149
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1644511149
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1644511149
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1644511149
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1644511149
transform 1 0 4048 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1644511149
transform 1 0 5152 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_57
timestamp 1644511149
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_69
timestamp 1644511149
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1644511149
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_113
timestamp 1644511149
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_125
timestamp 1644511149
transform 1 0 12604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_137
timestamp 1644511149
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_181
timestamp 1644511149
transform 1 0 17756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_193
timestamp 1644511149
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_200
timestamp 1644511149
transform 1 0 19504 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_212
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1644511149
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1644511149
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1644511149
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_281
timestamp 1644511149
transform 1 0 26956 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_293
timestamp 1644511149
transform 1 0 28060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_305
timestamp 1644511149
transform 1 0 29164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1644511149
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_393
timestamp 1644511149
transform 1 0 37260 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_405
timestamp 1644511149
transform 1 0 38364 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_417
timestamp 1644511149
transform 1 0 39468 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_439
timestamp 1644511149
transform 1 0 41492 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_447
timestamp 1644511149
transform 1 0 42228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_449
timestamp 1644511149
transform 1 0 42412 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_461
timestamp 1644511149
transform 1 0 43516 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1644511149
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_501
timestamp 1644511149
transform 1 0 47196 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_505
timestamp 1644511149
transform 1 0 47564 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_517
timestamp 1644511149
transform 1 0 48668 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_521
timestamp 1644511149
transform 1 0 49036 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_529
timestamp 1644511149
transform 1 0 49772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_533
timestamp 1644511149
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_545
timestamp 1644511149
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_557
timestamp 1644511149
transform 1 0 52348 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_561
timestamp 1644511149
transform 1 0 52716 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_573
timestamp 1644511149
transform 1 0 53820 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_585
timestamp 1644511149
transform 1 0 54924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_589
timestamp 1644511149
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_597
timestamp 1644511149
transform 1 0 56028 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_602
timestamp 1644511149
transform 1 0 56488 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_614
timestamp 1644511149
transform 1 0 57592 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1644511149
transform 1 0 57868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  Flash_110 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_111
timestamp 1644511149
transform 1 0 26220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_112
timestamp 1644511149
transform 1 0 41216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_113
timestamp 1644511149
transform 1 0 48760 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_114
timestamp 1644511149
transform 1 0 56212 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_115
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_116
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_117
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_118
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_119
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_120
timestamp 1644511149
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_121
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_122
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_123
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_124
timestamp 1644511149
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_125
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_126
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_127
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_128
timestamp 1644511149
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_129
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_130
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_131
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_132
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_133
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_134
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_135
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_136
timestamp 1644511149
transform 1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_137
timestamp 1644511149
transform 1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_138
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_139
timestamp 1644511149
transform 1 0 35328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_140
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_141
timestamp 1644511149
transform 1 0 38548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_142
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_143
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_144
timestamp 1644511149
transform 1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_145
timestamp 1644511149
transform 1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_146
timestamp 1644511149
transform 1 0 45816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_147
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_148
timestamp 1644511149
transform 1 0 48760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_149
timestamp 1644511149
transform 1 0 49956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_150
timestamp 1644511149
transform 1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_151
timestamp 1644511149
transform 1 0 52900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_152
timestamp 1644511149
transform 1 0 54372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_153
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_154
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_155
timestamp 1644511149
transform 1 0 57960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_156
timestamp 1644511149
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_157
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_158
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_159
timestamp 1644511149
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_160
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_161
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_162
timestamp 1644511149
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_163
timestamp 1644511149
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 16560 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 21712 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 26864 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 37168 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 42320 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 47472 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 52624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 57776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _220_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _221_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _222_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _223_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 1644511149
transform 1 0 15180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _226_
timestamp 1644511149
transform 1 0 12328 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _227_
timestamp 1644511149
transform 1 0 14260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _228_
timestamp 1644511149
transform 1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _229_
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _230_
timestamp 1644511149
transform 1 0 14996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _232_
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _233_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _234_
timestamp 1644511149
transform 1 0 9384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp 1644511149
transform 1 0 14444 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _236_
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _237_
timestamp 1644511149
transform 1 0 6532 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _238_
timestamp 1644511149
transform 1 0 17112 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _239_
timestamp 1644511149
transform 1 0 14076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _240_
timestamp 1644511149
transform 1 0 7728 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _241_
timestamp 1644511149
transform 1 0 7360 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _242_
timestamp 1644511149
transform 1 0 7452 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _243_
timestamp 1644511149
transform 1 0 12696 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _244_
timestamp 1644511149
transform 1 0 7084 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1644511149
transform 1 0 8004 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _246_
timestamp 1644511149
transform 1 0 14536 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _247_
timestamp 1644511149
transform 1 0 8004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _248_
timestamp 1644511149
transform 1 0 8280 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _249_
timestamp 1644511149
transform 1 0 13432 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _250_
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1644511149
transform 1 0 9568 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _253_
timestamp 1644511149
transform 1 0 7268 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _254_
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _255_
timestamp 1644511149
transform 1 0 18400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _256_
timestamp 1644511149
transform 1 0 7728 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _257_
timestamp 1644511149
transform 1 0 10212 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _258_
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _259_
timestamp 1644511149
transform 1 0 20332 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _261_
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _262_
timestamp 1644511149
transform 1 0 10304 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _263_
timestamp 1644511149
transform 1 0 19412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1644511149
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _265_
timestamp 1644511149
transform 1 0 7268 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _266_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _267_
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _268_
timestamp 1644511149
transform 1 0 6624 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _269_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1644511149
transform 1 0 7452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _271_
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _272_
timestamp 1644511149
transform 1 0 17664 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _273_
timestamp 1644511149
transform 1 0 9844 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _274_
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _275_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _276_
timestamp 1644511149
transform 1 0 10120 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _277_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _278_
timestamp 1644511149
transform 1 0 15640 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _279_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _280_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _281_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6808 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  _282_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1932 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _283_
timestamp 1644511149
transform 1 0 2944 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _284_
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _285_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _289_
timestamp 1644511149
transform 1 0 2576 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _291_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _292_
timestamp 1644511149
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _293_
timestamp 1644511149
transform 1 0 2208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1644511149
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1644511149
transform 1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _299_
timestamp 1644511149
transform 1 0 2300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1644511149
transform 1 0 5336 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1644511149
transform 1 0 5520 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp 1644511149
transform 1 0 4140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _304_
timestamp 1644511149
transform 1 0 2116 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1644511149
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp 1644511149
transform 1 0 2208 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _307_
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1644511149
transform 1 0 2208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1644511149
transform 1 0 2208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _310_
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp 1644511149
transform 1 0 2208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp 1644511149
transform 1 0 4600 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _314_
timestamp 1644511149
transform 1 0 3404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1644511149
transform 1 0 2208 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1644511149
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1644511149
transform 1 0 3404 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1644511149
transform 1 0 3680 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _319_
timestamp 1644511149
transform 1 0 2208 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp 1644511149
transform 1 0 2208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _321_
timestamp 1644511149
transform 1 0 3496 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp 1644511149
transform 1 0 3956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _323_
timestamp 1644511149
transform 1 0 2392 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _325_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _328_
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp 1644511149
transform 1 0 2852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1644511149
transform 1 0 4508 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1644511149
transform 1 0 4784 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1644511149
transform 1 0 2392 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1644511149
transform 1 0 2208 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _335_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _336_
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _337_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _338_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp 1644511149
transform 1 0 2668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _340_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _341_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp 1644511149
transform 1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp 1644511149
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1644511149
transform 1 0 12788 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1644511149
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1644511149
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _349_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _350_
timestamp 1644511149
transform 1 0 4508 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _351_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _353_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _355_
timestamp 1644511149
transform 1 0 7544 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _356_
timestamp 1644511149
transform 1 0 4968 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _357_
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _358_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _359_
timestamp 1644511149
transform 1 0 4232 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _360_
timestamp 1644511149
transform 1 0 4232 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1644511149
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _363_
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _365_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _367_
timestamp 1644511149
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _368_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _369_
timestamp 1644511149
transform 1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _370_
timestamp 1644511149
transform 1 0 8280 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _371_
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _372_
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _373_
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _374_
timestamp 1644511149
transform 1 0 8464 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _375_
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _376_
timestamp 1644511149
transform 1 0 9752 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _377_
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _378_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _379_
timestamp 1644511149
transform 1 0 10120 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _380_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _381_
timestamp 1644511149
transform 1 0 10028 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _382_
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _383_
timestamp 1644511149
transform 1 0 13156 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_2  _384_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _385_
timestamp 1644511149
transform 1 0 15824 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _386_
timestamp 1644511149
transform 1 0 14628 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _387_
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _388_
timestamp 1644511149
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _389_
timestamp 1644511149
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _390_
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _391_
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _392_
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _393_
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _394_
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _395_
timestamp 1644511149
transform 1 0 10488 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _396_
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _397_
timestamp 1644511149
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _398_
timestamp 1644511149
transform 1 0 10764 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _399_
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _400_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _401_
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _402_
timestamp 1644511149
transform 1 0 12696 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _403_
timestamp 1644511149
transform 1 0 10120 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _404_
timestamp 1644511149
transform 1 0 13064 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _405_
timestamp 1644511149
transform 1 0 12604 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _406_
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _407_
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _408_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _409_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _410_
timestamp 1644511149
transform 1 0 16744 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _411_
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _412_
timestamp 1644511149
transform 1 0 13248 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _413_
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _414_
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _415_
timestamp 1644511149
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _416_
timestamp 1644511149
transform 1 0 15272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _417_
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _418_
timestamp 1644511149
transform 1 0 15272 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _419_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _420_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _421_
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _422_
timestamp 1644511149
transform 1 0 17480 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _423_
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _424_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _425_
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _427_
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _428_
timestamp 1644511149
transform 1 0 16376 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _429_
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _430_
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _431_
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _432_
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _433_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _434_
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _435_
timestamp 1644511149
transform 1 0 17204 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _436_
timestamp 1644511149
transform 1 0 17204 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _437_
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _438_
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _439_
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _440_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _441_
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _442_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _443_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _444_
timestamp 1644511149
transform 1 0 14260 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _445_
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _446_
timestamp 1644511149
transform 1 0 14352 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _447_
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _448_
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _449_
timestamp 1644511149
transform 1 0 15456 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _450_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp 1644511149
transform 1 0 17020 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1644511149
transform 1 0 14536 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1644511149
transform 1 0 16836 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1644511149
transform 1 0 16652 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1644511149
transform 1 0 13432 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _465_
timestamp 1644511149
transform 1 0 15456 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _466_
timestamp 1644511149
transform 1 0 14352 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _467_
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _468_
timestamp 1644511149
transform 1 0 10948 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _469_
timestamp 1644511149
transform 1 0 9568 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _470_
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _471_
timestamp 1644511149
transform 1 0 6164 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _472_
timestamp 1644511149
transform 1 0 6992 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _473_
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _474_
timestamp 1644511149
transform 1 0 5888 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _475_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _476_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _477_
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _478_
timestamp 1644511149
transform 1 0 5244 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _479_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1644511149
transform 1 0 8740 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _481_
timestamp 1644511149
transform 1 0 12696 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _482_
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1644511149
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1644511149
transform 1 0 2392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1644511149
transform 1 0 1840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1644511149
transform 1 0 6256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1644511149
transform 1 0 4416 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1644511149
transform 1 0 5428 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1644511149
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1644511149
transform 1 0 1840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1644511149
transform 1 0 1932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1644511149
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1644511149
transform 1 0 1840 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1644511149
transform 1 0 4140 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1644511149
transform 1 0 1840 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1644511149
transform 1 0 3128 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1644511149
transform 1 0 2852 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1644511149
transform 1 0 6716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _508_
timestamp 1644511149
transform 1 0 3772 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1644511149
transform 1 0 6532 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1644511149
transform 1 0 17480 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1644511149
transform 1 0 13064 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _568_
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1644511149
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1644511149
transform 1 0 33396 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1644511149
transform 1 0 45080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1644511149
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1644511149
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1644511149
transform 1 0 50968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 53912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1644511149
transform 1 0 56764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1644511149
transform 1 0 56856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1644511149
transform 1 0 57684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 15916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 2852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input55 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 1656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 2852 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 2116 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3698 41200 3754 42000 6 flash_csb
port 0 nsew signal tristate
rlabel metal2 s 11150 41200 11206 42000 6 flash_io0_read
port 1 nsew signal input
rlabel metal2 s 18694 41200 18750 42000 6 flash_io0_we
port 2 nsew signal tristate
rlabel metal2 s 26146 41200 26202 42000 6 flash_io0_write
port 3 nsew signal tristate
rlabel metal2 s 33690 41200 33746 42000 6 flash_io1_read
port 4 nsew signal input
rlabel metal2 s 41142 41200 41198 42000 6 flash_io1_we
port 5 nsew signal tristate
rlabel metal2 s 48686 41200 48742 42000 6 flash_io1_write
port 6 nsew signal tristate
rlabel metal2 s 56138 41200 56194 42000 6 flash_sck
port 7 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 sram_addr0[0]
port 8 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 sram_addr0[1]
port 9 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 sram_addr0[2]
port 10 nsew signal tristate
rlabel metal2 s 11334 0 11390 800 6 sram_addr0[3]
port 11 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 sram_addr0[4]
port 12 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 sram_addr0[5]
port 13 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 sram_addr0[6]
port 14 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 sram_addr0[7]
port 15 nsew signal tristate
rlabel metal2 s 24030 0 24086 800 6 sram_addr0[8]
port 16 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 sram_addr1[0]
port 17 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 sram_addr1[1]
port 18 nsew signal tristate
rlabel metal2 s 8942 0 8998 800 6 sram_addr1[2]
port 19 nsew signal tristate
rlabel metal2 s 11886 0 11942 800 6 sram_addr1[3]
port 20 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 sram_addr1[4]
port 21 nsew signal tristate
rlabel metal2 s 17222 0 17278 800 6 sram_addr1[5]
port 22 nsew signal tristate
rlabel metal2 s 19706 0 19762 800 6 sram_addr1[6]
port 23 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 sram_addr1[7]
port 24 nsew signal tristate
rlabel metal2 s 24582 0 24638 800 6 sram_addr1[8]
port 25 nsew signal tristate
rlabel metal2 s 202 0 258 800 6 sram_clk0
port 26 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 sram_clk1
port 27 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 sram_csb0
port 28 nsew signal tristate
rlabel metal2 s 1582 0 1638 800 6 sram_csb1
port 29 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 sram_din0[0]
port 30 nsew signal tristate
rlabel metal2 s 27986 0 28042 800 6 sram_din0[10]
port 31 nsew signal tristate
rlabel metal2 s 29458 0 29514 800 6 sram_din0[11]
port 32 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 sram_din0[12]
port 33 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 sram_din0[13]
port 34 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 sram_din0[14]
port 35 nsew signal tristate
rlabel metal2 s 35254 0 35310 800 6 sram_din0[15]
port 36 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 sram_din0[16]
port 37 nsew signal tristate
rlabel metal2 s 38198 0 38254 800 6 sram_din0[17]
port 38 nsew signal tristate
rlabel metal2 s 39670 0 39726 800 6 sram_din0[18]
port 39 nsew signal tristate
rlabel metal2 s 41142 0 41198 800 6 sram_din0[19]
port 40 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 sram_din0[1]
port 41 nsew signal tristate
rlabel metal2 s 42614 0 42670 800 6 sram_din0[20]
port 42 nsew signal tristate
rlabel metal2 s 44086 0 44142 800 6 sram_din0[21]
port 43 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 sram_din0[22]
port 44 nsew signal tristate
rlabel metal2 s 46938 0 46994 800 6 sram_din0[23]
port 45 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 sram_din0[24]
port 46 nsew signal tristate
rlabel metal2 s 49882 0 49938 800 6 sram_din0[25]
port 47 nsew signal tristate
rlabel metal2 s 51354 0 51410 800 6 sram_din0[26]
port 48 nsew signal tristate
rlabel metal2 s 52826 0 52882 800 6 sram_din0[27]
port 49 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 sram_din0[28]
port 50 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 sram_din0[29]
port 51 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 sram_din0[2]
port 52 nsew signal tristate
rlabel metal2 s 57242 0 57298 800 6 sram_din0[30]
port 53 nsew signal tristate
rlabel metal2 s 58714 0 58770 800 6 sram_din0[31]
port 54 nsew signal tristate
rlabel metal2 s 12346 0 12402 800 6 sram_din0[3]
port 55 nsew signal tristate
rlabel metal2 s 15290 0 15346 800 6 sram_din0[4]
port 56 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 sram_din0[5]
port 57 nsew signal tristate
rlabel metal2 s 20166 0 20222 800 6 sram_din0[6]
port 58 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 sram_din0[7]
port 59 nsew signal tristate
rlabel metal2 s 25042 0 25098 800 6 sram_din0[8]
port 60 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 sram_din0[9]
port 61 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 sram_dout0[0]
port 62 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 sram_dout0[10]
port 63 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[11]
port 64 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 sram_dout0[12]
port 65 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sram_dout0[13]
port 66 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 sram_dout0[14]
port 67 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 sram_dout0[15]
port 68 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 sram_dout0[16]
port 69 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 sram_dout0[17]
port 70 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 sram_dout0[18]
port 71 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 sram_dout0[19]
port 72 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 sram_dout0[1]
port 73 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 sram_dout0[20]
port 74 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 sram_dout0[21]
port 75 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 sram_dout0[22]
port 76 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout0[23]
port 77 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 sram_dout0[24]
port 78 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 sram_dout0[25]
port 79 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 sram_dout0[26]
port 80 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 sram_dout0[27]
port 81 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout0[28]
port 82 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 sram_dout0[29]
port 83 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 sram_dout0[2]
port 84 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 sram_dout0[30]
port 85 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 sram_dout0[31]
port 86 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 sram_dout0[3]
port 87 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 sram_dout0[4]
port 88 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 sram_dout0[5]
port 89 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 sram_dout0[6]
port 90 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 sram_dout0[7]
port 91 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 sram_dout0[8]
port 92 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 sram_dout0[9]
port 93 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 sram_dout1[0]
port 94 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 sram_dout1[10]
port 95 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 sram_dout1[11]
port 96 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 sram_dout1[12]
port 97 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 sram_dout1[13]
port 98 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 sram_dout1[14]
port 99 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 sram_dout1[15]
port 100 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 sram_dout1[16]
port 101 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 sram_dout1[17]
port 102 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 sram_dout1[18]
port 103 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 sram_dout1[19]
port 104 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 sram_dout1[1]
port 105 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 sram_dout1[20]
port 106 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 sram_dout1[21]
port 107 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 sram_dout1[22]
port 108 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 sram_dout1[23]
port 109 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 sram_dout1[24]
port 110 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 sram_dout1[25]
port 111 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[26]
port 112 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 sram_dout1[27]
port 113 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 sram_dout1[28]
port 114 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 sram_dout1[29]
port 115 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 sram_dout1[2]
port 116 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 sram_dout1[30]
port 117 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 sram_dout1[31]
port 118 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 sram_dout1[3]
port 119 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 sram_dout1[4]
port 120 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 sram_dout1[5]
port 121 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 sram_dout1[6]
port 122 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 sram_dout1[7]
port 123 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout1[8]
port 124 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 sram_dout1[9]
port 125 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 sram_web0
port 126 nsew signal tristate
rlabel metal2 s 5078 0 5134 800 6 sram_wmask0[0]
port 127 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 sram_wmask0[1]
port 128 nsew signal tristate
rlabel metal2 s 10874 0 10930 800 6 sram_wmask0[2]
port 129 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 sram_wmask0[3]
port 130 nsew signal tristate
rlabel metal4 s 4208 2128 4528 39760 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 39760 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 39760 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 39760 6 vssd1
port 132 nsew ground bidirectional
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 133 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 wb_adr_i[0]
port 134 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wb_adr_i[10]
port 135 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[11]
port 136 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[12]
port 137 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[13]
port 138 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[14]
port 139 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 wb_adr_i[15]
port 140 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 wb_adr_i[16]
port 141 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 wb_adr_i[17]
port 142 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 wb_adr_i[18]
port 143 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_adr_i[19]
port 144 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wb_adr_i[1]
port 145 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_adr_i[20]
port 146 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_adr_i[21]
port 147 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 wb_adr_i[22]
port 148 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[23]
port 149 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 wb_adr_i[2]
port 150 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 wb_adr_i[3]
port 151 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 wb_adr_i[4]
port 152 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 wb_adr_i[5]
port 153 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 wb_adr_i[6]
port 154 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wb_adr_i[7]
port 155 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 wb_adr_i[8]
port 156 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wb_adr_i[9]
port 157 nsew signal input
rlabel metal3 s 0 552 800 672 6 wb_clk_i
port 158 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wb_cyc_i
port 159 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 wb_data_i[0]
port 160 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wb_data_i[10]
port 161 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[11]
port 162 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[12]
port 163 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[13]
port 164 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[14]
port 165 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 wb_data_i[15]
port 166 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_data_i[16]
port 167 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 wb_data_i[17]
port 168 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 wb_data_i[18]
port 169 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 wb_data_i[19]
port 170 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 wb_data_i[1]
port 171 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[20]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 wb_data_i[21]
port 173 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 wb_data_i[22]
port 174 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 wb_data_i[23]
port 175 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wb_data_i[24]
port 176 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 wb_data_i[25]
port 177 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 wb_data_i[26]
port 178 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 wb_data_i[27]
port 179 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 wb_data_i[28]
port 180 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 wb_data_i[29]
port 181 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 wb_data_i[2]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 wb_data_i[30]
port 183 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 wb_data_i[31]
port 184 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 wb_data_i[3]
port 185 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_data_i[4]
port 186 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_data_i[5]
port 187 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_data_i[6]
port 188 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 wb_data_i[7]
port 189 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wb_data_i[8]
port 190 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wb_data_i[9]
port 191 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 wb_data_o[0]
port 192 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 wb_data_o[10]
port 193 nsew signal tristate
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[11]
port 194 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[12]
port 195 nsew signal tristate
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[13]
port 196 nsew signal tristate
rlabel metal3 s 0 23672 800 23792 6 wb_data_o[14]
port 197 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 wb_data_o[15]
port 198 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wb_data_o[16]
port 199 nsew signal tristate
rlabel metal3 s 0 27344 800 27464 6 wb_data_o[17]
port 200 nsew signal tristate
rlabel metal3 s 0 28704 800 28824 6 wb_data_o[18]
port 201 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 wb_data_o[19]
port 202 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 wb_data_o[1]
port 203 nsew signal tristate
rlabel metal3 s 0 31152 800 31272 6 wb_data_o[20]
port 204 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[21]
port 205 nsew signal tristate
rlabel metal3 s 0 33736 800 33856 6 wb_data_o[22]
port 206 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wb_data_o[23]
port 207 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wb_data_o[24]
port 208 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wb_data_o[25]
port 209 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wb_data_o[26]
port 210 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wb_data_o[27]
port 211 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wb_data_o[28]
port 212 nsew signal tristate
rlabel metal3 s 0 39992 800 40112 6 wb_data_o[29]
port 213 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 wb_data_o[2]
port 214 nsew signal tristate
rlabel metal3 s 0 40808 800 40928 6 wb_data_o[30]
port 215 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 wb_data_o[31]
port 216 nsew signal tristate
rlabel metal3 s 0 9256 800 9376 6 wb_data_o[3]
port 217 nsew signal tristate
rlabel metal3 s 0 11024 800 11144 6 wb_data_o[4]
port 218 nsew signal tristate
rlabel metal3 s 0 12248 800 12368 6 wb_data_o[5]
port 219 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 wb_data_o[6]
port 220 nsew signal tristate
rlabel metal3 s 0 14832 800 14952 6 wb_data_o[7]
port 221 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 wb_data_o[8]
port 222 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 wb_data_o[9]
port 223 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wb_error_o
port 224 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 wb_rst_i
port 225 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 wb_sel_i[0]
port 226 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_sel_i[1]
port 227 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 wb_sel_i[2]
port 228 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_sel_i[3]
port 229 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wb_stall_o
port 230 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 wb_stb_i
port 231 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 42000
<< end >>
