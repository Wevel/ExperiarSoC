magic
tech sky130A
magscale 1 2
timestamp 1651190563
<< obsli1 >>
rect 1104 2159 78844 92497
<< obsm1 >>
rect 1104 2128 78844 92528
<< metal2 >>
rect 19982 0 20038 800
rect 60002 0 60058 800
<< obsm2 >>
rect 1308 856 78548 94217
rect 1308 711 19926 856
rect 20094 711 59946 856
rect 60114 711 78548 856
<< metal3 >>
rect 0 94120 800 94240
rect 79200 93440 80000 93560
rect 0 92488 800 92608
rect 0 90856 800 90976
rect 79200 90448 80000 90568
rect 0 89224 800 89344
rect 0 87592 800 87712
rect 79200 87456 80000 87576
rect 0 85960 800 86080
rect 0 84464 800 84584
rect 79200 84464 80000 84584
rect 0 82832 800 82952
rect 79200 81472 80000 81592
rect 0 81200 800 81320
rect 0 79568 800 79688
rect 79200 78480 80000 78600
rect 0 77936 800 78056
rect 0 76304 800 76424
rect 79200 75624 80000 75744
rect 0 74672 800 74792
rect 0 73176 800 73296
rect 79200 72632 80000 72752
rect 0 71544 800 71664
rect 0 69912 800 70032
rect 79200 69640 80000 69760
rect 0 68280 800 68400
rect 0 66648 800 66768
rect 79200 66648 80000 66768
rect 0 65016 800 65136
rect 0 63520 800 63640
rect 79200 63656 80000 63776
rect 0 61888 800 62008
rect 79200 60664 80000 60784
rect 0 60256 800 60376
rect 0 58624 800 58744
rect 79200 57808 80000 57928
rect 0 56992 800 57112
rect 0 55360 800 55480
rect 79200 54816 80000 54936
rect 0 53728 800 53848
rect 0 52232 800 52352
rect 79200 51824 80000 51944
rect 0 50600 800 50720
rect 0 48968 800 49088
rect 79200 48832 80000 48952
rect 0 47336 800 47456
rect 0 45704 800 45824
rect 79200 45840 80000 45960
rect 0 44072 800 44192
rect 79200 42848 80000 42968
rect 0 42576 800 42696
rect 0 40944 800 41064
rect 79200 39856 80000 39976
rect 0 39312 800 39432
rect 0 37680 800 37800
rect 79200 37000 80000 37120
rect 0 36048 800 36168
rect 0 34416 800 34536
rect 79200 34008 80000 34128
rect 0 32784 800 32904
rect 0 31288 800 31408
rect 79200 31016 80000 31136
rect 0 29656 800 29776
rect 0 28024 800 28144
rect 79200 28024 80000 28144
rect 0 26392 800 26512
rect 79200 25032 80000 25152
rect 0 24760 800 24880
rect 0 23128 800 23248
rect 79200 22040 80000 22160
rect 0 21632 800 21752
rect 0 20000 800 20120
rect 79200 19184 80000 19304
rect 0 18368 800 18488
rect 0 16736 800 16856
rect 79200 16192 80000 16312
rect 0 15104 800 15224
rect 0 13472 800 13592
rect 79200 13200 80000 13320
rect 0 11840 800 11960
rect 0 10344 800 10464
rect 79200 10208 80000 10328
rect 0 8712 800 8832
rect 0 7080 800 7200
rect 79200 7216 80000 7336
rect 0 5448 800 5568
rect 79200 4224 80000 4344
rect 0 3816 800 3936
rect 0 2184 800 2304
rect 79200 1368 80000 1488
rect 0 688 800 808
<< obsm3 >>
rect 880 94040 79200 94213
rect 800 93640 79200 94040
rect 800 93360 79120 93640
rect 800 92688 79200 93360
rect 880 92408 79200 92688
rect 800 91056 79200 92408
rect 880 90776 79200 91056
rect 800 90648 79200 90776
rect 800 90368 79120 90648
rect 800 89424 79200 90368
rect 880 89144 79200 89424
rect 800 87792 79200 89144
rect 880 87656 79200 87792
rect 880 87512 79120 87656
rect 800 87376 79120 87512
rect 800 86160 79200 87376
rect 880 85880 79200 86160
rect 800 84664 79200 85880
rect 880 84384 79120 84664
rect 800 83032 79200 84384
rect 880 82752 79200 83032
rect 800 81672 79200 82752
rect 800 81400 79120 81672
rect 880 81392 79120 81400
rect 880 81120 79200 81392
rect 800 79768 79200 81120
rect 880 79488 79200 79768
rect 800 78680 79200 79488
rect 800 78400 79120 78680
rect 800 78136 79200 78400
rect 880 77856 79200 78136
rect 800 76504 79200 77856
rect 880 76224 79200 76504
rect 800 75824 79200 76224
rect 800 75544 79120 75824
rect 800 74872 79200 75544
rect 880 74592 79200 74872
rect 800 73376 79200 74592
rect 880 73096 79200 73376
rect 800 72832 79200 73096
rect 800 72552 79120 72832
rect 800 71744 79200 72552
rect 880 71464 79200 71744
rect 800 70112 79200 71464
rect 880 69840 79200 70112
rect 880 69832 79120 69840
rect 800 69560 79120 69832
rect 800 68480 79200 69560
rect 880 68200 79200 68480
rect 800 66848 79200 68200
rect 880 66568 79120 66848
rect 800 65216 79200 66568
rect 880 64936 79200 65216
rect 800 63856 79200 64936
rect 800 63720 79120 63856
rect 880 63576 79120 63720
rect 880 63440 79200 63576
rect 800 62088 79200 63440
rect 880 61808 79200 62088
rect 800 60864 79200 61808
rect 800 60584 79120 60864
rect 800 60456 79200 60584
rect 880 60176 79200 60456
rect 800 58824 79200 60176
rect 880 58544 79200 58824
rect 800 58008 79200 58544
rect 800 57728 79120 58008
rect 800 57192 79200 57728
rect 880 56912 79200 57192
rect 800 55560 79200 56912
rect 880 55280 79200 55560
rect 800 55016 79200 55280
rect 800 54736 79120 55016
rect 800 53928 79200 54736
rect 880 53648 79200 53928
rect 800 52432 79200 53648
rect 880 52152 79200 52432
rect 800 52024 79200 52152
rect 800 51744 79120 52024
rect 800 50800 79200 51744
rect 880 50520 79200 50800
rect 800 49168 79200 50520
rect 880 49032 79200 49168
rect 880 48888 79120 49032
rect 800 48752 79120 48888
rect 800 47536 79200 48752
rect 880 47256 79200 47536
rect 800 46040 79200 47256
rect 800 45904 79120 46040
rect 880 45760 79120 45904
rect 880 45624 79200 45760
rect 800 44272 79200 45624
rect 880 43992 79200 44272
rect 800 43048 79200 43992
rect 800 42776 79120 43048
rect 880 42768 79120 42776
rect 880 42496 79200 42768
rect 800 41144 79200 42496
rect 880 40864 79200 41144
rect 800 40056 79200 40864
rect 800 39776 79120 40056
rect 800 39512 79200 39776
rect 880 39232 79200 39512
rect 800 37880 79200 39232
rect 880 37600 79200 37880
rect 800 37200 79200 37600
rect 800 36920 79120 37200
rect 800 36248 79200 36920
rect 880 35968 79200 36248
rect 800 34616 79200 35968
rect 880 34336 79200 34616
rect 800 34208 79200 34336
rect 800 33928 79120 34208
rect 800 32984 79200 33928
rect 880 32704 79200 32984
rect 800 31488 79200 32704
rect 880 31216 79200 31488
rect 880 31208 79120 31216
rect 800 30936 79120 31208
rect 800 29856 79200 30936
rect 880 29576 79200 29856
rect 800 28224 79200 29576
rect 880 27944 79120 28224
rect 800 26592 79200 27944
rect 880 26312 79200 26592
rect 800 25232 79200 26312
rect 800 24960 79120 25232
rect 880 24952 79120 24960
rect 880 24680 79200 24952
rect 800 23328 79200 24680
rect 880 23048 79200 23328
rect 800 22240 79200 23048
rect 800 21960 79120 22240
rect 800 21832 79200 21960
rect 880 21552 79200 21832
rect 800 20200 79200 21552
rect 880 19920 79200 20200
rect 800 19384 79200 19920
rect 800 19104 79120 19384
rect 800 18568 79200 19104
rect 880 18288 79200 18568
rect 800 16936 79200 18288
rect 880 16656 79200 16936
rect 800 16392 79200 16656
rect 800 16112 79120 16392
rect 800 15304 79200 16112
rect 880 15024 79200 15304
rect 800 13672 79200 15024
rect 880 13400 79200 13672
rect 880 13392 79120 13400
rect 800 13120 79120 13392
rect 800 12040 79200 13120
rect 880 11760 79200 12040
rect 800 10544 79200 11760
rect 880 10408 79200 10544
rect 880 10264 79120 10408
rect 800 10128 79120 10264
rect 800 8912 79200 10128
rect 880 8632 79200 8912
rect 800 7416 79200 8632
rect 800 7280 79120 7416
rect 880 7136 79120 7280
rect 880 7000 79200 7136
rect 800 5648 79200 7000
rect 880 5368 79200 5648
rect 800 4424 79200 5368
rect 800 4144 79120 4424
rect 800 4016 79200 4144
rect 880 3736 79200 4016
rect 800 2384 79200 3736
rect 880 2104 79200 2384
rect 800 1568 79200 2104
rect 800 1288 79120 1568
rect 800 888 79200 1288
rect 880 715 79200 888
<< metal4 >>
rect 4208 2128 4528 92528
rect 19568 2128 19888 92528
rect 34928 2128 35248 92528
rect 50288 2128 50608 92528
rect 65648 2128 65968 92528
<< obsm4 >>
rect 1715 2347 4128 89861
rect 4608 2347 19488 89861
rect 19968 2347 34848 89861
rect 35328 2347 50208 89861
rect 50688 2347 65568 89861
rect 66048 2347 77221 89861
<< labels >>
rlabel metal2 s 19982 0 20038 800 6 clk
port 1 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 peripheralBus_address[0]
port 2 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 peripheralBus_address[10]
port 3 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 peripheralBus_address[11]
port 4 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 peripheralBus_address[12]
port 5 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 peripheralBus_address[13]
port 6 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 peripheralBus_address[14]
port 7 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 peripheralBus_address[15]
port 8 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 peripheralBus_address[16]
port 9 nsew signal input
rlabel metal3 s 0 60256 800 60376 6 peripheralBus_address[17]
port 10 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 peripheralBus_address[18]
port 11 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 peripheralBus_address[19]
port 12 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 peripheralBus_address[1]
port 13 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 peripheralBus_address[20]
port 14 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 peripheralBus_address[21]
port 15 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 peripheralBus_address[22]
port 16 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 peripheralBus_address[23]
port 17 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 peripheralBus_address[2]
port 18 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 peripheralBus_address[3]
port 19 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 peripheralBus_address[4]
port 20 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 peripheralBus_address[5]
port 21 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 peripheralBus_address[6]
port 22 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 peripheralBus_address[7]
port 23 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 peripheralBus_address[8]
port 24 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 peripheralBus_address[9]
port 25 nsew signal input
rlabel metal3 s 0 688 800 808 6 peripheralBus_busy
port 26 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 peripheralBus_data[0]
port 27 nsew signal bidirectional
rlabel metal3 s 0 39312 800 39432 6 peripheralBus_data[10]
port 28 nsew signal bidirectional
rlabel metal3 s 0 42576 800 42696 6 peripheralBus_data[11]
port 29 nsew signal bidirectional
rlabel metal3 s 0 45704 800 45824 6 peripheralBus_data[12]
port 30 nsew signal bidirectional
rlabel metal3 s 0 48968 800 49088 6 peripheralBus_data[13]
port 31 nsew signal bidirectional
rlabel metal3 s 0 52232 800 52352 6 peripheralBus_data[14]
port 32 nsew signal bidirectional
rlabel metal3 s 0 55360 800 55480 6 peripheralBus_data[15]
port 33 nsew signal bidirectional
rlabel metal3 s 0 58624 800 58744 6 peripheralBus_data[16]
port 34 nsew signal bidirectional
rlabel metal3 s 0 61888 800 62008 6 peripheralBus_data[17]
port 35 nsew signal bidirectional
rlabel metal3 s 0 65016 800 65136 6 peripheralBus_data[18]
port 36 nsew signal bidirectional
rlabel metal3 s 0 68280 800 68400 6 peripheralBus_data[19]
port 37 nsew signal bidirectional
rlabel metal3 s 0 10344 800 10464 6 peripheralBus_data[1]
port 38 nsew signal bidirectional
rlabel metal3 s 0 71544 800 71664 6 peripheralBus_data[20]
port 39 nsew signal bidirectional
rlabel metal3 s 0 74672 800 74792 6 peripheralBus_data[21]
port 40 nsew signal bidirectional
rlabel metal3 s 0 77936 800 78056 6 peripheralBus_data[22]
port 41 nsew signal bidirectional
rlabel metal3 s 0 81200 800 81320 6 peripheralBus_data[23]
port 42 nsew signal bidirectional
rlabel metal3 s 0 82832 800 82952 6 peripheralBus_data[24]
port 43 nsew signal bidirectional
rlabel metal3 s 0 84464 800 84584 6 peripheralBus_data[25]
port 44 nsew signal bidirectional
rlabel metal3 s 0 85960 800 86080 6 peripheralBus_data[26]
port 45 nsew signal bidirectional
rlabel metal3 s 0 87592 800 87712 6 peripheralBus_data[27]
port 46 nsew signal bidirectional
rlabel metal3 s 0 89224 800 89344 6 peripheralBus_data[28]
port 47 nsew signal bidirectional
rlabel metal3 s 0 90856 800 90976 6 peripheralBus_data[29]
port 48 nsew signal bidirectional
rlabel metal3 s 0 13472 800 13592 6 peripheralBus_data[2]
port 49 nsew signal bidirectional
rlabel metal3 s 0 92488 800 92608 6 peripheralBus_data[30]
port 50 nsew signal bidirectional
rlabel metal3 s 0 94120 800 94240 6 peripheralBus_data[31]
port 51 nsew signal bidirectional
rlabel metal3 s 0 16736 800 16856 6 peripheralBus_data[3]
port 52 nsew signal bidirectional
rlabel metal3 s 0 20000 800 20120 6 peripheralBus_data[4]
port 53 nsew signal bidirectional
rlabel metal3 s 0 23128 800 23248 6 peripheralBus_data[5]
port 54 nsew signal bidirectional
rlabel metal3 s 0 26392 800 26512 6 peripheralBus_data[6]
port 55 nsew signal bidirectional
rlabel metal3 s 0 29656 800 29776 6 peripheralBus_data[7]
port 56 nsew signal bidirectional
rlabel metal3 s 0 32784 800 32904 6 peripheralBus_data[8]
port 57 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 peripheralBus_data[9]
port 58 nsew signal bidirectional
rlabel metal3 s 0 2184 800 2304 6 peripheralBus_oe
port 59 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 peripheralBus_we
port 60 nsew signal input
rlabel metal3 s 79200 1368 80000 1488 6 pwm_en[0]
port 61 nsew signal output
rlabel metal3 s 79200 60664 80000 60784 6 pwm_en[10]
port 62 nsew signal output
rlabel metal3 s 79200 66648 80000 66768 6 pwm_en[11]
port 63 nsew signal output
rlabel metal3 s 79200 72632 80000 72752 6 pwm_en[12]
port 64 nsew signal output
rlabel metal3 s 79200 78480 80000 78600 6 pwm_en[13]
port 65 nsew signal output
rlabel metal3 s 79200 84464 80000 84584 6 pwm_en[14]
port 66 nsew signal output
rlabel metal3 s 79200 90448 80000 90568 6 pwm_en[15]
port 67 nsew signal output
rlabel metal3 s 79200 7216 80000 7336 6 pwm_en[1]
port 68 nsew signal output
rlabel metal3 s 79200 13200 80000 13320 6 pwm_en[2]
port 69 nsew signal output
rlabel metal3 s 79200 19184 80000 19304 6 pwm_en[3]
port 70 nsew signal output
rlabel metal3 s 79200 25032 80000 25152 6 pwm_en[4]
port 71 nsew signal output
rlabel metal3 s 79200 31016 80000 31136 6 pwm_en[5]
port 72 nsew signal output
rlabel metal3 s 79200 37000 80000 37120 6 pwm_en[6]
port 73 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 pwm_en[7]
port 74 nsew signal output
rlabel metal3 s 79200 48832 80000 48952 6 pwm_en[8]
port 75 nsew signal output
rlabel metal3 s 79200 54816 80000 54936 6 pwm_en[9]
port 76 nsew signal output
rlabel metal3 s 79200 4224 80000 4344 6 pwm_out[0]
port 77 nsew signal output
rlabel metal3 s 79200 63656 80000 63776 6 pwm_out[10]
port 78 nsew signal output
rlabel metal3 s 79200 69640 80000 69760 6 pwm_out[11]
port 79 nsew signal output
rlabel metal3 s 79200 75624 80000 75744 6 pwm_out[12]
port 80 nsew signal output
rlabel metal3 s 79200 81472 80000 81592 6 pwm_out[13]
port 81 nsew signal output
rlabel metal3 s 79200 87456 80000 87576 6 pwm_out[14]
port 82 nsew signal output
rlabel metal3 s 79200 93440 80000 93560 6 pwm_out[15]
port 83 nsew signal output
rlabel metal3 s 79200 10208 80000 10328 6 pwm_out[1]
port 84 nsew signal output
rlabel metal3 s 79200 16192 80000 16312 6 pwm_out[2]
port 85 nsew signal output
rlabel metal3 s 79200 22040 80000 22160 6 pwm_out[3]
port 86 nsew signal output
rlabel metal3 s 79200 28024 80000 28144 6 pwm_out[4]
port 87 nsew signal output
rlabel metal3 s 79200 34008 80000 34128 6 pwm_out[5]
port 88 nsew signal output
rlabel metal3 s 79200 39856 80000 39976 6 pwm_out[6]
port 89 nsew signal output
rlabel metal3 s 79200 45840 80000 45960 6 pwm_out[7]
port 90 nsew signal output
rlabel metal3 s 79200 51824 80000 51944 6 pwm_out[8]
port 91 nsew signal output
rlabel metal3 s 79200 57808 80000 57928 6 pwm_out[9]
port 92 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 rst
port 93 nsew signal input
rlabel metal4 s 4208 2128 4528 92528 6 vccd1
port 94 nsew power input
rlabel metal4 s 34928 2128 35248 92528 6 vccd1
port 94 nsew power input
rlabel metal4 s 65648 2128 65968 92528 6 vccd1
port 94 nsew power input
rlabel metal4 s 19568 2128 19888 92528 6 vssd1
port 95 nsew ground input
rlabel metal4 s 50288 2128 50608 92528 6 vssd1
port 95 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 95000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22318100
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_PWM/runs/Peripheral_PWM/results/finishing/PWM.magic.gds
string GDS_START 580374
<< end >>

