magic
tech sky130A
magscale 1 2
timestamp 1653062880
<< viali >>
rect 1593 37417 1627 37451
rect 3433 37417 3467 37451
rect 14657 37417 14691 37451
rect 22937 37417 22971 37451
rect 27169 37417 27203 37451
rect 31217 37417 31251 37451
rect 35357 37417 35391 37451
rect 1961 37349 1995 37383
rect 2421 37349 2455 37383
rect 2789 37349 2823 37383
rect 3157 37349 3191 37383
rect 52009 37281 52043 37315
rect 76573 37281 76607 37315
rect 93409 37281 93443 37315
rect 1409 37213 1443 37247
rect 10333 37213 10367 37247
rect 39957 37213 39991 37247
rect 47593 37213 47627 37247
rect 51825 37213 51859 37247
rect 55873 37213 55907 37247
rect 60473 37213 60507 37247
rect 64153 37213 64187 37247
rect 68293 37213 68327 37247
rect 76849 37213 76883 37247
rect 84853 37213 84887 37247
rect 93225 37213 93259 37247
rect 109693 37213 109727 37247
rect 117881 37213 117915 37247
rect 40509 37145 40543 37179
rect 47777 37077 47811 37111
rect 56057 37077 56091 37111
rect 60657 37077 60691 37111
rect 64337 37077 64371 37111
rect 68477 37077 68511 37111
rect 85037 37077 85071 37111
rect 109877 37077 109911 37111
rect 117513 37077 117547 37111
rect 118065 37077 118099 37111
rect 1593 36873 1627 36907
rect 118065 36873 118099 36907
rect 1409 36737 1443 36771
rect 117513 36737 117547 36771
rect 117881 36737 117915 36771
rect 2053 36533 2087 36567
rect 2421 36533 2455 36567
rect 2789 36533 2823 36567
rect 3157 36533 3191 36567
rect 3525 36533 3559 36567
rect 1501 36125 1535 36159
rect 2053 36057 2087 36091
rect 117513 35037 117547 35071
rect 117881 35037 117915 35071
rect 118065 34901 118099 34935
rect 1409 34561 1443 34595
rect 1593 34357 1627 34391
rect 117881 33949 117915 33983
rect 117513 33813 117547 33847
rect 118065 33813 118099 33847
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 1409 29597 1443 29631
rect 117973 29529 118007 29563
rect 1593 29461 1627 29495
rect 118065 29461 118099 29495
rect 117881 26945 117915 26979
rect 117513 26741 117547 26775
rect 118065 26741 118099 26775
rect 1409 25857 1443 25891
rect 1685 25789 1719 25823
rect 1409 24157 1443 24191
rect 1593 24021 1627 24055
rect 117881 23681 117915 23715
rect 118065 23545 118099 23579
rect 117513 23477 117547 23511
rect 1409 22593 1443 22627
rect 117881 22593 117915 22627
rect 1685 22525 1719 22559
rect 117513 22389 117547 22423
rect 118065 22389 118099 22423
rect 117789 20825 117823 20859
rect 117881 20757 117915 20791
rect 68661 20553 68695 20587
rect 69213 20553 69247 20587
rect 70777 20553 70811 20587
rect 74181 20553 74215 20587
rect 74641 20553 74675 20587
rect 68569 20485 68603 20519
rect 65809 20417 65843 20451
rect 69653 20417 69687 20451
rect 73721 20417 73755 20451
rect 74549 20417 74583 20451
rect 65165 20349 65199 20383
rect 65901 20349 65935 20383
rect 66085 20349 66119 20383
rect 68753 20349 68787 20383
rect 69397 20349 69431 20383
rect 74733 20349 74767 20383
rect 65441 20213 65475 20247
rect 68201 20213 68235 20247
rect 73537 20213 73571 20247
rect 64981 20009 65015 20043
rect 68845 20009 68879 20043
rect 74917 20009 74951 20043
rect 73537 19873 73571 19907
rect 63601 19805 63635 19839
rect 69029 19805 69063 19839
rect 73793 19805 73827 19839
rect 63868 19737 63902 19771
rect 64245 19465 64279 19499
rect 66085 19465 66119 19499
rect 66821 19465 66855 19499
rect 69765 19465 69799 19499
rect 71145 19465 71179 19499
rect 118065 19465 118099 19499
rect 1685 19397 1719 19431
rect 68630 19397 68664 19431
rect 1409 19329 1443 19363
rect 64429 19329 64463 19363
rect 65993 19329 66027 19363
rect 67005 19329 67039 19363
rect 70685 19329 70719 19363
rect 70869 19329 70903 19363
rect 70961 19329 70995 19363
rect 117881 19329 117915 19363
rect 66177 19261 66211 19295
rect 68385 19261 68419 19295
rect 65625 19193 65659 19227
rect 70685 19125 70719 19159
rect 57345 18649 57379 18683
rect 57621 18581 57655 18615
rect 117789 18241 117823 18275
rect 117881 18037 117915 18071
rect 1409 17629 1443 17663
rect 1593 17493 1627 17527
rect 117789 15385 117823 15419
rect 117881 15317 117915 15351
rect 1869 14297 1903 14331
rect 1961 14229 1995 14263
rect 117237 12121 117271 12155
rect 117973 12121 118007 12155
rect 1869 11033 1903 11067
rect 2053 11033 2087 11067
rect 1409 9537 1443 9571
rect 1593 9333 1627 9367
rect 21833 8449 21867 8483
rect 22109 8381 22143 8415
rect 1593 7837 1627 7871
rect 1409 7701 1443 7735
rect 117973 6681 118007 6715
rect 118065 6613 118099 6647
rect 76665 6409 76699 6443
rect 77125 6409 77159 6443
rect 76021 6273 76055 6307
rect 77033 6273 77067 6307
rect 77217 6205 77251 6239
rect 75837 6069 75871 6103
rect 10057 5661 10091 5695
rect 17233 5661 17267 5695
rect 75929 5661 75963 5695
rect 76185 5661 76219 5695
rect 9873 5525 9907 5559
rect 17049 5525 17083 5559
rect 77309 5525 77343 5559
rect 9873 5321 9907 5355
rect 10333 5321 10367 5355
rect 17141 5321 17175 5355
rect 27905 5321 27939 5355
rect 28733 5321 28767 5355
rect 39221 5321 39255 5355
rect 39681 5321 39715 5355
rect 49985 5321 50019 5355
rect 50905 5321 50939 5355
rect 63969 5321 64003 5355
rect 64429 5321 64463 5355
rect 70041 5321 70075 5355
rect 70501 5321 70535 5355
rect 75837 5321 75871 5355
rect 92029 5321 92063 5355
rect 100677 5321 100711 5355
rect 17601 5253 17635 5287
rect 50813 5253 50847 5287
rect 76205 5253 76239 5287
rect 76297 5253 76331 5287
rect 10241 5185 10275 5219
rect 17509 5185 17543 5219
rect 21281 5185 21315 5219
rect 22201 5185 22235 5219
rect 28641 5185 28675 5219
rect 38761 5185 38795 5219
rect 39589 5185 39623 5219
rect 48872 5185 48906 5219
rect 53573 5185 53607 5219
rect 63233 5185 63267 5219
rect 64337 5185 64371 5219
rect 68753 5185 68787 5219
rect 70409 5185 70443 5219
rect 73629 5185 73663 5219
rect 75561 5185 75595 5219
rect 91937 5185 91971 5219
rect 96988 5185 97022 5219
rect 100769 5185 100803 5219
rect 102589 5185 102623 5219
rect 106729 5185 106763 5219
rect 117881 5185 117915 5219
rect 10517 5117 10551 5151
rect 17785 5117 17819 5151
rect 22293 5117 22327 5151
rect 22477 5117 22511 5151
rect 28917 5117 28951 5151
rect 39865 5117 39899 5151
rect 48605 5117 48639 5151
rect 50997 5117 51031 5151
rect 53757 5117 53791 5151
rect 64521 5117 64555 5151
rect 70593 5117 70627 5151
rect 76389 5117 76423 5151
rect 92121 5117 92155 5151
rect 96721 5117 96755 5151
rect 100309 5117 100343 5151
rect 100493 5117 100527 5151
rect 102333 5117 102367 5151
rect 106473 5117 106507 5151
rect 21833 5049 21867 5083
rect 22845 5049 22879 5083
rect 21097 4981 21131 5015
rect 28273 4981 28307 5015
rect 38577 4981 38611 5015
rect 50445 4981 50479 5015
rect 63049 4981 63083 5015
rect 68569 4981 68603 5015
rect 73445 4981 73479 5015
rect 91569 4981 91603 5015
rect 98101 4981 98135 5015
rect 103713 4981 103747 5015
rect 107853 4981 107887 5015
rect 118065 4981 118099 5015
rect 18429 4777 18463 4811
rect 22661 4777 22695 4811
rect 49341 4777 49375 4811
rect 63049 4777 63083 4811
rect 69213 4777 69247 4811
rect 76941 4777 76975 4811
rect 90833 4777 90867 4811
rect 97181 4777 97215 4811
rect 100217 4777 100251 4811
rect 104541 4777 104575 4811
rect 104909 4709 104943 4743
rect 27537 4641 27571 4675
rect 50169 4641 50203 4675
rect 52745 4641 52779 4675
rect 61669 4641 61703 4675
rect 76757 4641 76791 4675
rect 89453 4641 89487 4675
rect 97641 4641 97675 4675
rect 105001 4641 105035 4675
rect 112453 4641 112487 4675
rect 112545 4641 112579 4675
rect 9597 4573 9631 4607
rect 17049 4573 17083 4607
rect 17305 4573 17339 4607
rect 21281 4573 21315 4607
rect 21537 4573 21571 4607
rect 29745 4573 29779 4607
rect 49525 4573 49559 4607
rect 50353 4573 50387 4607
rect 52561 4573 52595 4607
rect 61936 4573 61970 4607
rect 67833 4573 67867 4607
rect 68100 4573 68134 4607
rect 72709 4573 72743 4607
rect 72976 4573 73010 4607
rect 76941 4573 76975 4607
rect 93961 4573 93995 4607
rect 94145 4573 94179 4607
rect 97365 4573 97399 4607
rect 97549 4573 97583 4607
rect 100217 4573 100251 4607
rect 100401 4573 100435 4607
rect 104725 4573 104759 4607
rect 107393 4573 107427 4607
rect 111349 4573 111383 4607
rect 9864 4505 9898 4539
rect 27804 4505 27838 4539
rect 76481 4505 76515 4539
rect 89720 4505 89754 4539
rect 94329 4505 94363 4539
rect 10977 4437 11011 4471
rect 28917 4437 28951 4471
rect 29561 4437 29595 4471
rect 50537 4437 50571 4471
rect 74089 4437 74123 4471
rect 77125 4437 77159 4471
rect 107209 4437 107243 4471
rect 111165 4437 111199 4471
rect 111993 4437 112027 4471
rect 112361 4437 112395 4471
rect 39957 4233 39991 4267
rect 86877 4233 86911 4267
rect 90373 4233 90407 4267
rect 100401 4233 100435 4267
rect 104357 4233 104391 4267
rect 112085 4233 112119 4267
rect 72433 4165 72467 4199
rect 97549 4165 97583 4199
rect 101321 4165 101355 4199
rect 107362 4165 107396 4199
rect 110972 4165 111006 4199
rect 117973 4165 118007 4199
rect 10241 4097 10275 4131
rect 10333 4097 10367 4131
rect 19717 4097 19751 4131
rect 19901 4097 19935 4131
rect 22937 4097 22971 4131
rect 28365 4097 28399 4131
rect 38833 4097 38867 4131
rect 63233 4097 63267 4131
rect 68385 4097 68419 4131
rect 72801 4097 72835 4131
rect 73905 4097 73939 4131
rect 73997 4097 74031 4131
rect 77309 4097 77343 4131
rect 86233 4097 86267 4131
rect 87245 4097 87279 4131
rect 90557 4097 90591 4131
rect 91201 4097 91235 4131
rect 94053 4097 94087 4131
rect 97273 4097 97307 4131
rect 100217 4097 100251 4131
rect 100493 4097 100527 4131
rect 100953 4097 100987 4131
rect 101137 4097 101171 4131
rect 101505 4097 101539 4131
rect 101781 4097 101815 4131
rect 104265 4097 104299 4131
rect 104449 4097 104483 4131
rect 104909 4097 104943 4131
rect 105093 4097 105127 4131
rect 118157 4097 118191 4131
rect 22753 4029 22787 4063
rect 28181 4029 28215 4063
rect 38577 4029 38611 4063
rect 63049 4029 63083 4063
rect 68201 4029 68235 4063
rect 77585 4029 77619 4063
rect 86509 4029 86543 4063
rect 87337 4029 87371 4063
rect 87521 4029 87555 4063
rect 94329 4029 94363 4063
rect 100033 4029 100067 4063
rect 107117 4029 107151 4063
rect 110705 4029 110739 4063
rect 10517 3893 10551 3927
rect 20085 3893 20119 3927
rect 23121 3893 23155 3927
rect 28549 3893 28583 3927
rect 63417 3893 63451 3927
rect 68569 3893 68603 3927
rect 74181 3893 74215 3927
rect 86049 3893 86083 3927
rect 89361 3893 89395 3927
rect 91017 3893 91051 3927
rect 104909 3893 104943 3927
rect 108497 3893 108531 3927
rect 59277 3689 59311 3723
rect 83749 3689 83783 3723
rect 91753 3689 91787 3723
rect 92489 3689 92523 3723
rect 98009 3689 98043 3723
rect 100125 3689 100159 3723
rect 107301 3689 107335 3723
rect 112269 3689 112303 3723
rect 45661 3621 45695 3655
rect 46489 3621 46523 3655
rect 92213 3621 92247 3655
rect 94329 3621 94363 3655
rect 99113 3621 99147 3655
rect 52745 3553 52779 3587
rect 54125 3553 54159 3587
rect 56149 3553 56183 3587
rect 64337 3553 64371 3587
rect 83657 3553 83691 3587
rect 86233 3553 86267 3587
rect 91937 3553 91971 3587
rect 93961 3553 93995 3587
rect 97181 3553 97215 3587
rect 101689 3553 101723 3587
rect 102174 3553 102208 3587
rect 107853 3553 107887 3587
rect 112361 3553 112395 3587
rect 1409 3485 1443 3519
rect 2421 3485 2455 3519
rect 10149 3485 10183 3519
rect 19993 3485 20027 3519
rect 23765 3485 23799 3519
rect 28549 3485 28583 3519
rect 38485 3485 38519 3519
rect 38597 3485 38631 3519
rect 45477 3485 45511 3519
rect 46305 3485 46339 3519
rect 47409 3485 47443 3519
rect 47593 3485 47627 3519
rect 50169 3485 50203 3519
rect 52469 3485 52503 3519
rect 55965 3485 55999 3519
rect 59093 3485 59127 3519
rect 62221 3485 62255 3519
rect 64061 3485 64095 3519
rect 66085 3485 66119 3519
rect 67833 3485 67867 3519
rect 74181 3485 74215 3519
rect 83565 3485 83599 3519
rect 86489 3485 86523 3519
rect 88717 3485 88751 3519
rect 89085 3485 89119 3519
rect 89453 3485 89487 3519
rect 90005 3485 90039 3519
rect 92069 3485 92103 3519
rect 95157 3485 95191 3519
rect 97089 3485 97123 3519
rect 100125 3485 100159 3519
rect 100309 3485 100343 3519
rect 102057 3485 102091 3519
rect 107669 3485 107703 3519
rect 108681 3485 108715 3519
rect 112140 3485 112174 3519
rect 117881 3485 117915 3519
rect 2881 3417 2915 3451
rect 37657 3417 37691 3451
rect 37841 3417 37875 3451
rect 47777 3417 47811 3451
rect 53389 3417 53423 3451
rect 66453 3417 66487 3451
rect 68201 3417 68235 3451
rect 90649 3417 90683 3451
rect 91569 3417 91603 3451
rect 91753 3417 91787 3451
rect 92397 3417 92431 3451
rect 97917 3417 97951 3451
rect 98837 3417 98871 3451
rect 111993 3417 112027 3451
rect 1593 3349 1627 3383
rect 2237 3349 2271 3383
rect 9965 3349 9999 3383
rect 19809 3349 19843 3383
rect 23581 3349 23615 3383
rect 28365 3349 28399 3383
rect 38761 3349 38795 3383
rect 50353 3349 50387 3383
rect 62313 3349 62347 3383
rect 73997 3349 74031 3383
rect 83933 3349 83967 3383
rect 87613 3349 87647 3383
rect 94421 3349 94455 3383
rect 94973 3349 95007 3383
rect 96629 3349 96663 3383
rect 96997 3349 97031 3383
rect 101965 3349 101999 3383
rect 102333 3349 102367 3383
rect 107761 3349 107795 3383
rect 108497 3349 108531 3383
rect 112637 3349 112671 3383
rect 118065 3349 118099 3383
rect 2237 3145 2271 3179
rect 52009 3145 52043 3179
rect 53297 3145 53331 3179
rect 54953 3145 54987 3179
rect 57897 3145 57931 3179
rect 66361 3145 66395 3179
rect 68385 3145 68419 3179
rect 113373 3145 113407 3179
rect 118065 3145 118099 3179
rect 56977 3077 57011 3111
rect 83933 3077 83967 3111
rect 94228 3077 94262 3111
rect 100861 3077 100895 3111
rect 111800 3077 111834 3111
rect 1409 3009 1443 3043
rect 2421 3009 2455 3043
rect 2881 3009 2915 3043
rect 22201 3009 22235 3043
rect 28457 3009 28491 3043
rect 32321 3009 32355 3043
rect 34989 3009 35023 3043
rect 40049 3009 40083 3043
rect 43361 3009 43395 3043
rect 47777 3009 47811 3043
rect 50261 3009 50295 3043
rect 50629 3009 50663 3043
rect 52193 3009 52227 3043
rect 52929 3009 52963 3043
rect 53113 3009 53147 3043
rect 54769 3009 54803 3043
rect 55965 3009 55999 3043
rect 56701 3009 56735 3043
rect 56793 3009 56827 3043
rect 58081 3009 58115 3043
rect 59829 3009 59863 3043
rect 61117 3009 61151 3043
rect 63233 3009 63267 3043
rect 66269 3009 66303 3043
rect 68201 3009 68235 3043
rect 69305 3009 69339 3043
rect 70593 3009 70627 3043
rect 73629 3009 73663 3043
rect 74365 3009 74399 3043
rect 76573 3009 76607 3043
rect 79701 3009 79735 3043
rect 83657 3009 83691 3043
rect 86233 3009 86267 3043
rect 86601 3009 86635 3043
rect 86877 3009 86911 3043
rect 87429 3009 87463 3043
rect 89361 3009 89395 3043
rect 89545 3009 89579 3043
rect 90189 3009 90223 3043
rect 91201 3009 91235 3043
rect 92029 3009 92063 3043
rect 93961 3009 93995 3043
rect 97089 3009 97123 3043
rect 99573 3009 99607 3043
rect 100125 3009 100159 3043
rect 100769 3009 100803 3043
rect 104265 3009 104299 3043
rect 105185 3009 105219 3043
rect 107301 3009 107335 3043
rect 107568 3009 107602 3043
rect 111073 3009 111107 3043
rect 113557 3009 113591 3043
rect 114845 3009 114879 3043
rect 117973 3009 118007 3043
rect 8401 2941 8435 2975
rect 32137 2941 32171 2975
rect 39865 2941 39899 2975
rect 43177 2941 43211 2975
rect 44189 2941 44223 2975
rect 47593 2941 47627 2975
rect 47961 2941 47995 2975
rect 55781 2941 55815 2975
rect 56149 2941 56183 2975
rect 61853 2941 61887 2975
rect 69581 2941 69615 2975
rect 70777 2941 70811 2975
rect 79977 2941 80011 2975
rect 87613 2941 87647 2975
rect 88993 2941 89027 2975
rect 89177 2941 89211 2975
rect 101045 2941 101079 2975
rect 111533 2941 111567 2975
rect 43545 2873 43579 2907
rect 73813 2873 73847 2907
rect 86049 2873 86083 2907
rect 91017 2873 91051 2907
rect 97273 2873 97307 2907
rect 108681 2873 108715 2907
rect 110889 2873 110923 2907
rect 1593 2805 1627 2839
rect 3065 2805 3099 2839
rect 22017 2805 22051 2839
rect 28641 2805 28675 2839
rect 29377 2805 29411 2839
rect 31585 2805 31619 2839
rect 32505 2805 32539 2839
rect 34805 2805 34839 2839
rect 35817 2805 35851 2839
rect 37473 2805 37507 2839
rect 39773 2805 39807 2839
rect 40233 2805 40267 2839
rect 51273 2805 51307 2839
rect 59645 2805 59679 2839
rect 63049 2805 63083 2839
rect 65441 2805 65475 2839
rect 74549 2805 74583 2839
rect 75285 2805 75319 2839
rect 76389 2805 76423 2839
rect 77401 2805 77435 2839
rect 82185 2805 82219 2839
rect 90281 2805 90315 2839
rect 92121 2805 92155 2839
rect 95341 2805 95375 2839
rect 96629 2805 96663 2839
rect 99757 2805 99791 2839
rect 100401 2805 100435 2839
rect 104449 2805 104483 2839
rect 105369 2805 105403 2839
rect 112913 2805 112947 2839
rect 115029 2805 115063 2839
rect 22385 2601 22419 2635
rect 43729 2601 43763 2635
rect 49433 2601 49467 2635
rect 53113 2601 53147 2635
rect 85405 2601 85439 2635
rect 88165 2601 88199 2635
rect 89453 2601 89487 2635
rect 91753 2601 91787 2635
rect 93225 2601 93259 2635
rect 96905 2601 96939 2635
rect 108313 2601 108347 2635
rect 111073 2601 111107 2635
rect 33977 2533 34011 2567
rect 42717 2533 42751 2567
rect 61945 2533 61979 2567
rect 63417 2533 63451 2567
rect 65993 2533 66027 2567
rect 67281 2533 67315 2567
rect 69489 2533 69523 2567
rect 69949 2533 69983 2567
rect 71605 2533 71639 2567
rect 73721 2533 73755 2567
rect 83105 2533 83139 2567
rect 97733 2533 97767 2567
rect 98193 2533 98227 2567
rect 101873 2533 101907 2567
rect 106013 2533 106047 2567
rect 113373 2533 113407 2567
rect 2421 2465 2455 2499
rect 43361 2465 43395 2499
rect 63049 2465 63083 2499
rect 66453 2465 66487 2499
rect 66821 2465 66855 2499
rect 68845 2465 68879 2499
rect 70961 2465 70995 2499
rect 73353 2465 73387 2499
rect 74549 2465 74583 2499
rect 77033 2465 77067 2499
rect 92581 2465 92615 2499
rect 94789 2465 94823 2499
rect 97365 2465 97399 2499
rect 99113 2465 99147 2499
rect 104633 2465 104667 2499
rect 109969 2465 110003 2499
rect 111625 2465 111659 2499
rect 1409 2397 1443 2431
rect 4629 2397 4663 2431
rect 4997 2397 5031 2431
rect 5273 2397 5307 2431
rect 6561 2397 6595 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 11713 2397 11747 2431
rect 13921 2397 13955 2431
rect 14565 2397 14599 2431
rect 14841 2397 14875 2431
rect 15853 2397 15887 2431
rect 17417 2397 17451 2431
rect 18705 2397 18739 2431
rect 19625 2397 19659 2431
rect 20637 2397 20671 2431
rect 22017 2397 22051 2431
rect 22201 2397 22235 2431
rect 23857 2397 23891 2431
rect 24409 2397 24443 2431
rect 25421 2397 25455 2431
rect 27169 2397 27203 2431
rect 27813 2397 27847 2431
rect 28457 2397 28491 2431
rect 28641 2397 28675 2431
rect 28825 2397 28859 2431
rect 29561 2397 29595 2431
rect 31033 2397 31067 2431
rect 31401 2397 31435 2431
rect 31677 2397 31711 2431
rect 32873 2397 32907 2431
rect 34989 2397 35023 2431
rect 35173 2397 35207 2431
rect 35357 2397 35391 2431
rect 36277 2397 36311 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40417 2397 40451 2431
rect 40693 2397 40727 2431
rect 41613 2397 41647 2431
rect 42901 2397 42935 2431
rect 43545 2397 43579 2431
rect 44373 2397 44407 2431
rect 45385 2397 45419 2431
rect 46213 2397 46247 2431
rect 47041 2397 47075 2431
rect 47593 2397 47627 2431
rect 47777 2397 47811 2431
rect 48605 2397 48639 2431
rect 49617 2397 49651 2431
rect 50997 2397 51031 2431
rect 52193 2397 52227 2431
rect 52745 2397 52779 2431
rect 52929 2397 52963 2431
rect 53757 2397 53791 2431
rect 54769 2397 54803 2431
rect 55781 2397 55815 2431
rect 56425 2397 56459 2431
rect 56609 2397 56643 2431
rect 58173 2397 58207 2431
rect 60657 2397 60691 2431
rect 61669 2397 61703 2431
rect 61761 2397 61795 2431
rect 63233 2397 63267 2431
rect 64061 2397 64095 2431
rect 64705 2397 64739 2431
rect 65625 2397 65659 2431
rect 65809 2397 65843 2431
rect 66637 2397 66671 2431
rect 67465 2397 67499 2431
rect 68569 2397 68603 2431
rect 68661 2397 68695 2431
rect 70133 2397 70167 2431
rect 71789 2397 71823 2431
rect 72617 2397 72651 2431
rect 73537 2397 73571 2431
rect 74733 2397 74767 2431
rect 74917 2397 74951 2431
rect 75929 2397 75963 2431
rect 77217 2397 77251 2431
rect 77401 2397 77435 2431
rect 78505 2397 78539 2431
rect 79425 2397 79459 2431
rect 80069 2397 80103 2431
rect 81449 2397 81483 2431
rect 81909 2397 81943 2431
rect 82093 2397 82127 2431
rect 82737 2397 82771 2431
rect 82921 2397 82955 2431
rect 83841 2397 83875 2431
rect 84577 2397 84611 2431
rect 86693 2397 86727 2431
rect 87889 2397 87923 2431
rect 87981 2397 88015 2431
rect 88993 2397 89027 2431
rect 89637 2397 89671 2431
rect 90557 2397 90591 2431
rect 90649 2397 90683 2431
rect 91385 2397 91419 2431
rect 91569 2397 91603 2431
rect 92305 2397 92339 2431
rect 92397 2397 92431 2431
rect 94145 2397 94179 2431
rect 95801 2397 95835 2431
rect 96537 2397 96571 2431
rect 96721 2397 96755 2431
rect 97549 2397 97583 2431
rect 98377 2397 98411 2431
rect 100953 2397 100987 2431
rect 101689 2397 101723 2431
rect 102241 2397 102275 2431
rect 102793 2397 102827 2431
rect 103345 2397 103379 2431
rect 104900 2397 104934 2431
rect 107577 2397 107611 2431
rect 108497 2397 108531 2431
rect 109785 2397 109819 2431
rect 110797 2397 110831 2431
rect 111441 2397 111475 2431
rect 112177 2397 112211 2431
rect 113189 2397 113223 2431
rect 114569 2397 114603 2431
rect 115581 2397 115615 2431
rect 115857 2397 115891 2431
rect 117145 2397 117179 2431
rect 117881 2397 117915 2431
rect 7757 2329 7791 2363
rect 12541 2329 12575 2363
rect 12725 2329 12759 2363
rect 29193 2329 29227 2363
rect 29837 2329 29871 2363
rect 33149 2329 33183 2363
rect 36001 2329 36035 2363
rect 36553 2329 36587 2363
rect 37933 2329 37967 2363
rect 39129 2329 39163 2363
rect 47961 2329 47995 2363
rect 50629 2329 50663 2363
rect 56793 2329 56827 2363
rect 59553 2329 59587 2363
rect 82277 2329 82311 2363
rect 85313 2329 85347 2363
rect 99380 2329 99414 2363
rect 103805 2329 103839 2363
rect 104449 2329 104483 2363
rect 3801 2261 3835 2295
rect 5457 2261 5491 2295
rect 7849 2261 7883 2295
rect 10241 2261 10275 2295
rect 13277 2261 13311 2295
rect 15025 2261 15059 2295
rect 17233 2261 17267 2295
rect 17877 2261 17911 2295
rect 19809 2261 19843 2295
rect 22845 2261 22879 2295
rect 24593 2261 24627 2295
rect 26985 2261 27019 2295
rect 30389 2261 30423 2295
rect 30665 2261 30699 2295
rect 30849 2261 30883 2295
rect 31861 2261 31895 2295
rect 32597 2261 32631 2295
rect 33701 2261 33735 2295
rect 37473 2261 37507 2295
rect 38393 2261 38427 2295
rect 39221 2261 39255 2295
rect 40877 2261 40911 2295
rect 44189 2261 44223 2295
rect 45201 2261 45235 2295
rect 46857 2261 46891 2295
rect 52009 2261 52043 2295
rect 54585 2261 54619 2295
rect 59829 2261 59863 2295
rect 64521 2261 64555 2295
rect 76113 2261 76147 2295
rect 78689 2261 78723 2295
rect 79241 2261 79275 2295
rect 81265 2261 81299 2295
rect 83657 2261 83691 2295
rect 86785 2261 86819 2295
rect 90833 2261 90867 2295
rect 93961 2261 93995 2295
rect 95617 2261 95651 2295
rect 100493 2261 100527 2295
rect 100769 2261 100803 2295
rect 101229 2261 101263 2295
rect 102977 2261 103011 2295
rect 107761 2261 107795 2295
rect 109417 2261 109451 2295
rect 109877 2261 109911 2295
rect 110613 2261 110647 2295
rect 111533 2261 111567 2295
rect 111993 2261 112027 2295
rect 112821 2261 112855 2295
rect 114753 2261 114787 2295
rect 117329 2261 117363 2295
rect 118065 2261 118099 2295
<< metal1 >>
rect 1104 37562 118864 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 96374 37562
rect 96426 37510 96438 37562
rect 96490 37510 96502 37562
rect 96554 37510 96566 37562
rect 96618 37510 96630 37562
rect 96682 37510 118864 37562
rect 1104 37488 118864 37510
rect 1578 37448 1584 37460
rect 1539 37420 1584 37448
rect 1578 37408 1584 37420
rect 1636 37408 1642 37460
rect 2038 37408 2044 37460
rect 2096 37448 2102 37460
rect 3421 37451 3479 37457
rect 3421 37448 3433 37451
rect 2096 37420 3433 37448
rect 2096 37408 2102 37420
rect 3421 37417 3433 37420
rect 3467 37417 3479 37451
rect 3421 37411 3479 37417
rect 14366 37408 14372 37460
rect 14424 37448 14430 37460
rect 14645 37451 14703 37457
rect 14645 37448 14657 37451
rect 14424 37420 14657 37448
rect 14424 37408 14430 37420
rect 14645 37417 14657 37420
rect 14691 37417 14703 37451
rect 14645 37411 14703 37417
rect 22646 37408 22652 37460
rect 22704 37448 22710 37460
rect 22925 37451 22983 37457
rect 22925 37448 22937 37451
rect 22704 37420 22937 37448
rect 22704 37408 22710 37420
rect 22925 37417 22937 37420
rect 22971 37417 22983 37451
rect 22925 37411 22983 37417
rect 26786 37408 26792 37460
rect 26844 37448 26850 37460
rect 27157 37451 27215 37457
rect 27157 37448 27169 37451
rect 26844 37420 27169 37448
rect 26844 37408 26850 37420
rect 27157 37417 27169 37420
rect 27203 37417 27215 37451
rect 27157 37411 27215 37417
rect 30926 37408 30932 37460
rect 30984 37448 30990 37460
rect 31205 37451 31263 37457
rect 31205 37448 31217 37451
rect 30984 37420 31217 37448
rect 30984 37408 30990 37420
rect 31205 37417 31217 37420
rect 31251 37417 31263 37451
rect 35342 37448 35348 37460
rect 35303 37420 35348 37448
rect 31205 37411 31263 37417
rect 35342 37408 35348 37420
rect 35400 37408 35406 37460
rect 1949 37383 2007 37389
rect 1949 37349 1961 37383
rect 1995 37380 2007 37383
rect 2409 37383 2467 37389
rect 2409 37380 2421 37383
rect 1995 37352 2421 37380
rect 1995 37349 2007 37352
rect 1949 37343 2007 37349
rect 2409 37349 2421 37352
rect 2455 37380 2467 37383
rect 2777 37383 2835 37389
rect 2777 37380 2789 37383
rect 2455 37352 2789 37380
rect 2455 37349 2467 37352
rect 2409 37343 2467 37349
rect 2777 37349 2789 37352
rect 2823 37380 2835 37383
rect 3145 37383 3203 37389
rect 3145 37380 3157 37383
rect 2823 37352 3157 37380
rect 2823 37349 2835 37352
rect 2777 37343 2835 37349
rect 3145 37349 3157 37352
rect 3191 37380 3203 37383
rect 86862 37380 86868 37392
rect 3191 37352 86868 37380
rect 3191 37349 3203 37352
rect 3145 37343 3203 37349
rect 1397 37247 1455 37253
rect 1397 37213 1409 37247
rect 1443 37244 1455 37247
rect 1964 37244 1992 37343
rect 86862 37340 86868 37352
rect 86920 37340 86926 37392
rect 50890 37272 50896 37324
rect 50948 37312 50954 37324
rect 51997 37315 52055 37321
rect 51997 37312 52009 37315
rect 50948 37284 52009 37312
rect 50948 37272 50954 37284
rect 51997 37281 52009 37284
rect 52043 37281 52055 37315
rect 51997 37275 52055 37281
rect 76466 37272 76472 37324
rect 76524 37312 76530 37324
rect 76561 37315 76619 37321
rect 76561 37312 76573 37315
rect 76524 37284 76573 37312
rect 76524 37272 76530 37284
rect 76561 37281 76573 37284
rect 76607 37281 76619 37315
rect 76561 37275 76619 37281
rect 92014 37272 92020 37324
rect 92072 37312 92078 37324
rect 93397 37315 93455 37321
rect 93397 37312 93409 37315
rect 92072 37284 93409 37312
rect 92072 37272 92078 37284
rect 93397 37281 93409 37284
rect 93443 37281 93455 37315
rect 93397 37275 93455 37281
rect 1443 37216 1992 37244
rect 1443 37213 1455 37216
rect 1397 37207 1455 37213
rect 10226 37204 10232 37256
rect 10284 37244 10290 37256
rect 10321 37247 10379 37253
rect 10321 37244 10333 37247
rect 10284 37216 10333 37244
rect 10284 37204 10290 37216
rect 10321 37213 10333 37216
rect 10367 37213 10379 37247
rect 10321 37207 10379 37213
rect 39206 37204 39212 37256
rect 39264 37244 39270 37256
rect 39945 37247 40003 37253
rect 39945 37244 39957 37247
rect 39264 37216 39957 37244
rect 39264 37204 39270 37216
rect 39945 37213 39957 37216
rect 39991 37213 40003 37247
rect 47578 37244 47584 37256
rect 47539 37216 47584 37244
rect 39945 37207 40003 37213
rect 47578 37204 47584 37216
rect 47636 37204 47642 37256
rect 51626 37204 51632 37256
rect 51684 37244 51690 37256
rect 51813 37247 51871 37253
rect 51813 37244 51825 37247
rect 51684 37216 51825 37244
rect 51684 37204 51690 37216
rect 51813 37213 51825 37216
rect 51859 37213 51871 37247
rect 51813 37207 51871 37213
rect 54938 37204 54944 37256
rect 54996 37244 55002 37256
rect 55861 37247 55919 37253
rect 55861 37244 55873 37247
rect 54996 37216 55873 37244
rect 54996 37204 55002 37216
rect 55861 37213 55873 37216
rect 55907 37213 55919 37247
rect 55861 37207 55919 37213
rect 59262 37204 59268 37256
rect 59320 37244 59326 37256
rect 60461 37247 60519 37253
rect 60461 37244 60473 37247
rect 59320 37216 60473 37244
rect 59320 37204 59326 37216
rect 60461 37213 60473 37216
rect 60507 37213 60519 37247
rect 64138 37244 64144 37256
rect 64099 37216 64144 37244
rect 60461 37207 60519 37213
rect 64138 37204 64144 37216
rect 64196 37204 64202 37256
rect 68186 37204 68192 37256
rect 68244 37244 68250 37256
rect 68281 37247 68339 37253
rect 68281 37244 68293 37247
rect 68244 37216 68293 37244
rect 68244 37204 68250 37216
rect 68281 37213 68293 37216
rect 68327 37213 68339 37247
rect 68281 37207 68339 37213
rect 74626 37204 74632 37256
rect 74684 37244 74690 37256
rect 76837 37247 76895 37253
rect 76837 37244 76849 37247
rect 74684 37216 76849 37244
rect 74684 37204 74690 37216
rect 76837 37213 76849 37216
rect 76883 37213 76895 37247
rect 84838 37244 84844 37256
rect 84799 37216 84844 37244
rect 76837 37207 76895 37213
rect 84838 37204 84844 37216
rect 84896 37204 84902 37256
rect 93026 37204 93032 37256
rect 93084 37244 93090 37256
rect 93213 37247 93271 37253
rect 93213 37244 93225 37247
rect 93084 37216 93225 37244
rect 93084 37204 93090 37216
rect 93213 37213 93225 37216
rect 93259 37213 93271 37247
rect 109678 37244 109684 37256
rect 109639 37216 109684 37244
rect 93213 37207 93271 37213
rect 109678 37204 109684 37216
rect 109736 37204 109742 37256
rect 117869 37247 117927 37253
rect 117869 37244 117881 37247
rect 117516 37216 117881 37244
rect 40494 37176 40500 37188
rect 40455 37148 40500 37176
rect 40494 37136 40500 37148
rect 40552 37136 40558 37188
rect 117516 37120 117544 37216
rect 117869 37213 117881 37216
rect 117915 37213 117927 37247
rect 117869 37207 117927 37213
rect 47486 37068 47492 37120
rect 47544 37108 47550 37120
rect 47765 37111 47823 37117
rect 47765 37108 47777 37111
rect 47544 37080 47777 37108
rect 47544 37068 47550 37080
rect 47765 37077 47777 37080
rect 47811 37077 47823 37111
rect 47765 37071 47823 37077
rect 55766 37068 55772 37120
rect 55824 37108 55830 37120
rect 56045 37111 56103 37117
rect 56045 37108 56057 37111
rect 55824 37080 56057 37108
rect 55824 37068 55830 37080
rect 56045 37077 56057 37080
rect 56091 37077 56103 37111
rect 56045 37071 56103 37077
rect 59906 37068 59912 37120
rect 59964 37108 59970 37120
rect 60645 37111 60703 37117
rect 60645 37108 60657 37111
rect 59964 37080 60657 37108
rect 59964 37068 59970 37080
rect 60645 37077 60657 37080
rect 60691 37077 60703 37111
rect 60645 37071 60703 37077
rect 64046 37068 64052 37120
rect 64104 37108 64110 37120
rect 64325 37111 64383 37117
rect 64325 37108 64337 37111
rect 64104 37080 64337 37108
rect 64104 37068 64110 37080
rect 64325 37077 64337 37080
rect 64371 37077 64383 37111
rect 64325 37071 64383 37077
rect 64414 37068 64420 37120
rect 64472 37108 64478 37120
rect 68465 37111 68523 37117
rect 68465 37108 68477 37111
rect 64472 37080 68477 37108
rect 64472 37068 64478 37080
rect 68465 37077 68477 37080
rect 68511 37077 68523 37111
rect 68465 37071 68523 37077
rect 84746 37068 84752 37120
rect 84804 37108 84810 37120
rect 85025 37111 85083 37117
rect 85025 37108 85037 37111
rect 84804 37080 85037 37108
rect 84804 37068 84810 37080
rect 85025 37077 85037 37080
rect 85071 37077 85083 37111
rect 85025 37071 85083 37077
rect 109586 37068 109592 37120
rect 109644 37108 109650 37120
rect 109865 37111 109923 37117
rect 109865 37108 109877 37111
rect 109644 37080 109877 37108
rect 109644 37068 109650 37080
rect 109865 37077 109877 37080
rect 109911 37077 109923 37111
rect 117498 37108 117504 37120
rect 117459 37080 117504 37108
rect 109865 37071 109923 37077
rect 117498 37068 117504 37080
rect 117556 37068 117562 37120
rect 117866 37068 117872 37120
rect 117924 37108 117930 37120
rect 118053 37111 118111 37117
rect 118053 37108 118065 37111
rect 117924 37080 118065 37108
rect 117924 37068 117930 37080
rect 118053 37077 118065 37080
rect 118099 37077 118111 37111
rect 118053 37071 118111 37077
rect 1104 37018 118864 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 81014 37018
rect 81066 36966 81078 37018
rect 81130 36966 81142 37018
rect 81194 36966 81206 37018
rect 81258 36966 81270 37018
rect 81322 36966 111734 37018
rect 111786 36966 111798 37018
rect 111850 36966 111862 37018
rect 111914 36966 111926 37018
rect 111978 36966 111990 37018
rect 112042 36966 118864 37018
rect 1104 36944 118864 36966
rect 1581 36907 1639 36913
rect 1581 36873 1593 36907
rect 1627 36904 1639 36907
rect 2774 36904 2780 36916
rect 1627 36876 2780 36904
rect 1627 36873 1639 36876
rect 1581 36867 1639 36873
rect 2774 36864 2780 36876
rect 2832 36864 2838 36916
rect 45554 36864 45560 36916
rect 45612 36904 45618 36916
rect 64138 36904 64144 36916
rect 45612 36876 64144 36904
rect 45612 36864 45618 36876
rect 64138 36864 64144 36876
rect 64196 36864 64202 36916
rect 66346 36864 66352 36916
rect 66404 36904 66410 36916
rect 84838 36904 84844 36916
rect 66404 36876 84844 36904
rect 66404 36864 66410 36876
rect 84838 36864 84844 36876
rect 84896 36864 84902 36916
rect 117222 36864 117228 36916
rect 117280 36904 117286 36916
rect 118053 36907 118111 36913
rect 118053 36904 118065 36907
rect 117280 36876 118065 36904
rect 117280 36864 117286 36876
rect 118053 36873 118065 36876
rect 118099 36873 118111 36907
rect 118053 36867 118111 36873
rect 40494 36796 40500 36848
rect 40552 36836 40558 36848
rect 101766 36836 101772 36848
rect 40552 36808 101772 36836
rect 40552 36796 40558 36808
rect 101766 36796 101772 36808
rect 101824 36796 101830 36848
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1443 36740 2084 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 2056 36573 2084 36740
rect 92106 36728 92112 36780
rect 92164 36768 92170 36780
rect 117501 36771 117559 36777
rect 117501 36768 117513 36771
rect 92164 36740 117513 36768
rect 92164 36728 92170 36740
rect 117501 36737 117513 36740
rect 117547 36768 117559 36771
rect 117869 36771 117927 36777
rect 117869 36768 117881 36771
rect 117547 36740 117881 36768
rect 117547 36737 117559 36740
rect 117501 36731 117559 36737
rect 117869 36737 117881 36740
rect 117915 36737 117927 36771
rect 117869 36731 117927 36737
rect 2041 36567 2099 36573
rect 2041 36533 2053 36567
rect 2087 36564 2099 36567
rect 2409 36567 2467 36573
rect 2409 36564 2421 36567
rect 2087 36536 2421 36564
rect 2087 36533 2099 36536
rect 2041 36527 2099 36533
rect 2409 36533 2421 36536
rect 2455 36564 2467 36567
rect 2777 36567 2835 36573
rect 2777 36564 2789 36567
rect 2455 36536 2789 36564
rect 2455 36533 2467 36536
rect 2409 36527 2467 36533
rect 2777 36533 2789 36536
rect 2823 36564 2835 36567
rect 3145 36567 3203 36573
rect 3145 36564 3157 36567
rect 2823 36536 3157 36564
rect 2823 36533 2835 36536
rect 2777 36527 2835 36533
rect 3145 36533 3157 36536
rect 3191 36564 3203 36567
rect 3513 36567 3571 36573
rect 3513 36564 3525 36567
rect 3191 36536 3525 36564
rect 3191 36533 3203 36536
rect 3145 36527 3203 36533
rect 3513 36533 3525 36536
rect 3559 36564 3571 36567
rect 88702 36564 88708 36576
rect 3559 36536 88708 36564
rect 3559 36533 3571 36536
rect 3513 36527 3571 36533
rect 88702 36524 88708 36536
rect 88760 36524 88766 36576
rect 1104 36474 118864 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 96374 36474
rect 96426 36422 96438 36474
rect 96490 36422 96502 36474
rect 96554 36422 96566 36474
rect 96618 36422 96630 36474
rect 96682 36422 118864 36474
rect 1104 36400 118864 36422
rect 1486 36156 1492 36168
rect 1447 36128 1492 36156
rect 1486 36116 1492 36128
rect 1544 36116 1550 36168
rect 2041 36091 2099 36097
rect 2041 36057 2053 36091
rect 2087 36088 2099 36091
rect 86494 36088 86500 36100
rect 2087 36060 86500 36088
rect 2087 36057 2099 36060
rect 2041 36051 2099 36057
rect 86494 36048 86500 36060
rect 86552 36048 86558 36100
rect 1104 35930 118864 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 81014 35930
rect 81066 35878 81078 35930
rect 81130 35878 81142 35930
rect 81194 35878 81206 35930
rect 81258 35878 81270 35930
rect 81322 35878 111734 35930
rect 111786 35878 111798 35930
rect 111850 35878 111862 35930
rect 111914 35878 111926 35930
rect 111978 35878 111990 35930
rect 112042 35878 118864 35930
rect 1104 35856 118864 35878
rect 1104 35386 118864 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 96374 35386
rect 96426 35334 96438 35386
rect 96490 35334 96502 35386
rect 96554 35334 96566 35386
rect 96618 35334 96630 35386
rect 96682 35334 118864 35386
rect 1104 35312 118864 35334
rect 90266 35028 90272 35080
rect 90324 35068 90330 35080
rect 117501 35071 117559 35077
rect 117501 35068 117513 35071
rect 90324 35040 117513 35068
rect 90324 35028 90330 35040
rect 117501 35037 117513 35040
rect 117547 35068 117559 35071
rect 117869 35071 117927 35077
rect 117869 35068 117881 35071
rect 117547 35040 117881 35068
rect 117547 35037 117559 35040
rect 117501 35031 117559 35037
rect 117869 35037 117881 35040
rect 117915 35037 117927 35071
rect 117869 35031 117927 35037
rect 118050 34932 118056 34944
rect 118011 34904 118056 34932
rect 118050 34892 118056 34904
rect 118108 34892 118114 34944
rect 1104 34842 118864 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 81014 34842
rect 81066 34790 81078 34842
rect 81130 34790 81142 34842
rect 81194 34790 81206 34842
rect 81258 34790 81270 34842
rect 81322 34790 111734 34842
rect 111786 34790 111798 34842
rect 111850 34790 111862 34842
rect 111914 34790 111926 34842
rect 111978 34790 111990 34842
rect 112042 34790 118864 34842
rect 1104 34768 118864 34790
rect 1394 34592 1400 34604
rect 1355 34564 1400 34592
rect 1394 34552 1400 34564
rect 1452 34552 1458 34604
rect 1578 34388 1584 34400
rect 1539 34360 1584 34388
rect 1578 34348 1584 34360
rect 1636 34348 1642 34400
rect 1104 34298 118864 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 96374 34298
rect 96426 34246 96438 34298
rect 96490 34246 96502 34298
rect 96554 34246 96566 34298
rect 96618 34246 96630 34298
rect 96682 34246 118864 34298
rect 1104 34224 118864 34246
rect 117869 33983 117927 33989
rect 117869 33980 117881 33983
rect 117516 33952 117881 33980
rect 92474 33804 92480 33856
rect 92532 33844 92538 33856
rect 117516 33853 117544 33952
rect 117869 33949 117881 33952
rect 117915 33949 117927 33983
rect 117869 33943 117927 33949
rect 117501 33847 117559 33853
rect 117501 33844 117513 33847
rect 92532 33816 117513 33844
rect 92532 33804 92538 33816
rect 117501 33813 117513 33816
rect 117547 33813 117559 33847
rect 118050 33844 118056 33856
rect 118011 33816 118056 33844
rect 117501 33807 117559 33813
rect 118050 33804 118056 33816
rect 118108 33804 118114 33856
rect 1104 33754 118864 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 81014 33754
rect 81066 33702 81078 33754
rect 81130 33702 81142 33754
rect 81194 33702 81206 33754
rect 81258 33702 81270 33754
rect 81322 33702 111734 33754
rect 111786 33702 111798 33754
rect 111850 33702 111862 33754
rect 111914 33702 111926 33754
rect 111978 33702 111990 33754
rect 112042 33702 118864 33754
rect 1104 33680 118864 33702
rect 1104 33210 118864 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 96374 33210
rect 96426 33158 96438 33210
rect 96490 33158 96502 33210
rect 96554 33158 96566 33210
rect 96618 33158 96630 33210
rect 96682 33158 118864 33210
rect 1104 33136 118864 33158
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 1486 32892 1492 32904
rect 1443 32864 1492 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 1486 32852 1492 32864
rect 1544 32852 1550 32904
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 1104 32666 118864 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 81014 32666
rect 81066 32614 81078 32666
rect 81130 32614 81142 32666
rect 81194 32614 81206 32666
rect 81258 32614 81270 32666
rect 81322 32614 111734 32666
rect 111786 32614 111798 32666
rect 111850 32614 111862 32666
rect 111914 32614 111926 32666
rect 111978 32614 111990 32666
rect 112042 32614 118864 32666
rect 1104 32592 118864 32614
rect 1104 32122 118864 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 96374 32122
rect 96426 32070 96438 32122
rect 96490 32070 96502 32122
rect 96554 32070 96566 32122
rect 96618 32070 96630 32122
rect 96682 32070 118864 32122
rect 1104 32048 118864 32070
rect 1104 31578 118864 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 81014 31578
rect 81066 31526 81078 31578
rect 81130 31526 81142 31578
rect 81194 31526 81206 31578
rect 81258 31526 81270 31578
rect 81322 31526 111734 31578
rect 111786 31526 111798 31578
rect 111850 31526 111862 31578
rect 111914 31526 111926 31578
rect 111978 31526 111990 31578
rect 112042 31526 118864 31578
rect 1104 31504 118864 31526
rect 1104 31034 118864 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 96374 31034
rect 96426 30982 96438 31034
rect 96490 30982 96502 31034
rect 96554 30982 96566 31034
rect 96618 30982 96630 31034
rect 96682 30982 118864 31034
rect 1104 30960 118864 30982
rect 1104 30490 118864 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 81014 30490
rect 81066 30438 81078 30490
rect 81130 30438 81142 30490
rect 81194 30438 81206 30490
rect 81258 30438 81270 30490
rect 81322 30438 111734 30490
rect 111786 30438 111798 30490
rect 111850 30438 111862 30490
rect 111914 30438 111926 30490
rect 111978 30438 111990 30490
rect 112042 30438 118864 30490
rect 1104 30416 118864 30438
rect 1104 29946 118864 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 96374 29946
rect 96426 29894 96438 29946
rect 96490 29894 96502 29946
rect 96554 29894 96566 29946
rect 96618 29894 96630 29946
rect 96682 29894 118864 29946
rect 1104 29872 118864 29894
rect 1397 29631 1455 29637
rect 1397 29597 1409 29631
rect 1443 29628 1455 29631
rect 2038 29628 2044 29640
rect 1443 29600 2044 29628
rect 1443 29597 1455 29600
rect 1397 29591 1455 29597
rect 2038 29588 2044 29600
rect 2096 29588 2102 29640
rect 117958 29560 117964 29572
rect 117919 29532 117964 29560
rect 117958 29520 117964 29532
rect 118016 29520 118022 29572
rect 1578 29492 1584 29504
rect 1539 29464 1584 29492
rect 1578 29452 1584 29464
rect 1636 29452 1642 29504
rect 112438 29452 112444 29504
rect 112496 29492 112502 29504
rect 118053 29495 118111 29501
rect 118053 29492 118065 29495
rect 112496 29464 118065 29492
rect 112496 29452 112502 29464
rect 118053 29461 118065 29464
rect 118099 29461 118111 29495
rect 118053 29455 118111 29461
rect 1104 29402 118864 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 81014 29402
rect 81066 29350 81078 29402
rect 81130 29350 81142 29402
rect 81194 29350 81206 29402
rect 81258 29350 81270 29402
rect 81322 29350 111734 29402
rect 111786 29350 111798 29402
rect 111850 29350 111862 29402
rect 111914 29350 111926 29402
rect 111978 29350 111990 29402
rect 112042 29350 118864 29402
rect 1104 29328 118864 29350
rect 1104 28858 118864 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 96374 28858
rect 96426 28806 96438 28858
rect 96490 28806 96502 28858
rect 96554 28806 96566 28858
rect 96618 28806 96630 28858
rect 96682 28806 118864 28858
rect 1104 28784 118864 28806
rect 1104 28314 118864 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 81014 28314
rect 81066 28262 81078 28314
rect 81130 28262 81142 28314
rect 81194 28262 81206 28314
rect 81258 28262 81270 28314
rect 81322 28262 111734 28314
rect 111786 28262 111798 28314
rect 111850 28262 111862 28314
rect 111914 28262 111926 28314
rect 111978 28262 111990 28314
rect 112042 28262 118864 28314
rect 1104 28240 118864 28262
rect 1104 27770 118864 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 96374 27770
rect 96426 27718 96438 27770
rect 96490 27718 96502 27770
rect 96554 27718 96566 27770
rect 96618 27718 96630 27770
rect 96682 27718 118864 27770
rect 1104 27696 118864 27718
rect 1104 27226 118864 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 81014 27226
rect 81066 27174 81078 27226
rect 81130 27174 81142 27226
rect 81194 27174 81206 27226
rect 81258 27174 81270 27226
rect 81322 27174 111734 27226
rect 111786 27174 111798 27226
rect 111850 27174 111862 27226
rect 111914 27174 111926 27226
rect 111978 27174 111990 27226
rect 112042 27174 118864 27226
rect 1104 27152 118864 27174
rect 117869 26979 117927 26985
rect 117869 26976 117881 26979
rect 117516 26948 117881 26976
rect 64322 26732 64328 26784
rect 64380 26772 64386 26784
rect 117516 26781 117544 26948
rect 117869 26945 117881 26948
rect 117915 26945 117927 26979
rect 117869 26939 117927 26945
rect 117501 26775 117559 26781
rect 117501 26772 117513 26775
rect 64380 26744 117513 26772
rect 64380 26732 64386 26744
rect 117501 26741 117513 26744
rect 117547 26741 117559 26775
rect 118050 26772 118056 26784
rect 118011 26744 118056 26772
rect 117501 26735 117559 26741
rect 118050 26732 118056 26744
rect 118108 26732 118114 26784
rect 1104 26682 118864 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 96374 26682
rect 96426 26630 96438 26682
rect 96490 26630 96502 26682
rect 96554 26630 96566 26682
rect 96618 26630 96630 26682
rect 96682 26630 118864 26682
rect 1104 26608 118864 26630
rect 1104 26138 118864 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 81014 26138
rect 81066 26086 81078 26138
rect 81130 26086 81142 26138
rect 81194 26086 81206 26138
rect 81258 26086 81270 26138
rect 81322 26086 111734 26138
rect 111786 26086 111798 26138
rect 111850 26086 111862 26138
rect 111914 26086 111926 26138
rect 111978 26086 111990 26138
rect 112042 26086 118864 26138
rect 1104 26064 118864 26086
rect 1394 25984 1400 26036
rect 1452 26024 1458 26036
rect 1762 26024 1768 26036
rect 1452 25996 1768 26024
rect 1452 25984 1458 25996
rect 1762 25984 1768 25996
rect 1820 25984 1826 26036
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 1670 25820 1676 25832
rect 1631 25792 1676 25820
rect 1670 25780 1676 25792
rect 1728 25780 1734 25832
rect 1104 25594 118864 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 96374 25594
rect 96426 25542 96438 25594
rect 96490 25542 96502 25594
rect 96554 25542 96566 25594
rect 96618 25542 96630 25594
rect 96682 25542 118864 25594
rect 1104 25520 118864 25542
rect 1104 25050 118864 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 81014 25050
rect 81066 24998 81078 25050
rect 81130 24998 81142 25050
rect 81194 24998 81206 25050
rect 81258 24998 81270 25050
rect 81322 24998 111734 25050
rect 111786 24998 111798 25050
rect 111850 24998 111862 25050
rect 111914 24998 111926 25050
rect 111978 24998 111990 25050
rect 112042 24998 118864 25050
rect 1104 24976 118864 24998
rect 1104 24506 118864 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 96374 24506
rect 96426 24454 96438 24506
rect 96490 24454 96502 24506
rect 96554 24454 96566 24506
rect 96618 24454 96630 24506
rect 96682 24454 118864 24506
rect 1104 24432 118864 24454
rect 1397 24191 1455 24197
rect 1397 24157 1409 24191
rect 1443 24188 1455 24191
rect 1854 24188 1860 24200
rect 1443 24160 1860 24188
rect 1443 24157 1455 24160
rect 1397 24151 1455 24157
rect 1854 24148 1860 24160
rect 1912 24148 1918 24200
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 1104 23962 118864 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 81014 23962
rect 81066 23910 81078 23962
rect 81130 23910 81142 23962
rect 81194 23910 81206 23962
rect 81258 23910 81270 23962
rect 81322 23910 111734 23962
rect 111786 23910 111798 23962
rect 111850 23910 111862 23962
rect 111914 23910 111926 23962
rect 111978 23910 111990 23962
rect 112042 23910 118864 23962
rect 1104 23888 118864 23910
rect 117869 23715 117927 23721
rect 117869 23712 117881 23715
rect 117516 23684 117881 23712
rect 54110 23468 54116 23520
rect 54168 23508 54174 23520
rect 117516 23517 117544 23684
rect 117869 23681 117881 23684
rect 117915 23681 117927 23715
rect 117869 23675 117927 23681
rect 118050 23576 118056 23588
rect 118011 23548 118056 23576
rect 118050 23536 118056 23548
rect 118108 23536 118114 23588
rect 117501 23511 117559 23517
rect 117501 23508 117513 23511
rect 54168 23480 117513 23508
rect 54168 23468 54174 23480
rect 117501 23477 117513 23480
rect 117547 23477 117559 23511
rect 117501 23471 117559 23477
rect 1104 23418 118864 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 96374 23418
rect 96426 23366 96438 23418
rect 96490 23366 96502 23418
rect 96554 23366 96566 23418
rect 96618 23366 96630 23418
rect 96682 23366 118864 23418
rect 1104 23344 118864 23366
rect 1104 22874 118864 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 81014 22874
rect 81066 22822 81078 22874
rect 81130 22822 81142 22874
rect 81194 22822 81206 22874
rect 81258 22822 81270 22874
rect 81322 22822 111734 22874
rect 111786 22822 111798 22874
rect 111850 22822 111862 22874
rect 111914 22822 111926 22874
rect 111978 22822 111990 22874
rect 112042 22822 118864 22874
rect 1104 22800 118864 22822
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 117869 22627 117927 22633
rect 117869 22624 117881 22627
rect 117516 22596 117881 22624
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 68646 22556 68652 22568
rect 1719 22528 68652 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 68646 22516 68652 22528
rect 68704 22516 68710 22568
rect 52730 22380 52736 22432
rect 52788 22420 52794 22432
rect 117516 22429 117544 22596
rect 117869 22593 117881 22596
rect 117915 22593 117927 22627
rect 117869 22587 117927 22593
rect 117501 22423 117559 22429
rect 117501 22420 117513 22423
rect 52788 22392 117513 22420
rect 52788 22380 52794 22392
rect 117501 22389 117513 22392
rect 117547 22389 117559 22423
rect 118050 22420 118056 22432
rect 118011 22392 118056 22420
rect 117501 22383 117559 22389
rect 118050 22380 118056 22392
rect 118108 22380 118114 22432
rect 1104 22330 118864 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 96374 22330
rect 96426 22278 96438 22330
rect 96490 22278 96502 22330
rect 96554 22278 96566 22330
rect 96618 22278 96630 22330
rect 96682 22278 118864 22330
rect 1104 22256 118864 22278
rect 1104 21786 118864 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 81014 21786
rect 81066 21734 81078 21786
rect 81130 21734 81142 21786
rect 81194 21734 81206 21786
rect 81258 21734 81270 21786
rect 81322 21734 111734 21786
rect 111786 21734 111798 21786
rect 111850 21734 111862 21786
rect 111914 21734 111926 21786
rect 111978 21734 111990 21786
rect 112042 21734 118864 21786
rect 1104 21712 118864 21734
rect 1104 21242 118864 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 96374 21242
rect 96426 21190 96438 21242
rect 96490 21190 96502 21242
rect 96554 21190 96566 21242
rect 96618 21190 96630 21242
rect 96682 21190 118864 21242
rect 1104 21168 118864 21190
rect 117774 20856 117780 20868
rect 117735 20828 117780 20856
rect 117774 20816 117780 20828
rect 117832 20816 117838 20868
rect 77110 20748 77116 20800
rect 77168 20788 77174 20800
rect 117869 20791 117927 20797
rect 117869 20788 117881 20791
rect 77168 20760 117881 20788
rect 77168 20748 77174 20760
rect 117869 20757 117881 20760
rect 117915 20757 117927 20791
rect 117869 20751 117927 20757
rect 1104 20698 118864 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 81014 20698
rect 81066 20646 81078 20698
rect 81130 20646 81142 20698
rect 81194 20646 81206 20698
rect 81258 20646 81270 20698
rect 81322 20646 111734 20698
rect 111786 20646 111798 20698
rect 111850 20646 111862 20698
rect 111914 20646 111926 20698
rect 111978 20646 111990 20698
rect 112042 20646 118864 20698
rect 1104 20624 118864 20646
rect 68646 20584 68652 20596
rect 68607 20556 68652 20584
rect 68646 20544 68652 20556
rect 68704 20584 68710 20596
rect 69201 20587 69259 20593
rect 69201 20584 69213 20587
rect 68704 20556 69213 20584
rect 68704 20544 68710 20556
rect 69201 20553 69213 20556
rect 69247 20553 69259 20587
rect 69201 20547 69259 20553
rect 69290 20544 69296 20596
rect 69348 20584 69354 20596
rect 70394 20584 70400 20596
rect 69348 20556 70400 20584
rect 69348 20544 69354 20556
rect 70394 20544 70400 20556
rect 70452 20544 70458 20596
rect 70765 20587 70823 20593
rect 70765 20553 70777 20587
rect 70811 20553 70823 20587
rect 70765 20547 70823 20553
rect 74169 20587 74227 20593
rect 74169 20553 74181 20587
rect 74215 20553 74227 20587
rect 74626 20584 74632 20596
rect 74587 20556 74632 20584
rect 74169 20547 74227 20553
rect 68557 20519 68615 20525
rect 68557 20485 68569 20519
rect 68603 20516 68615 20519
rect 70670 20516 70676 20528
rect 68603 20488 70676 20516
rect 68603 20485 68615 20488
rect 68557 20479 68615 20485
rect 70670 20476 70676 20488
rect 70728 20516 70734 20528
rect 70780 20516 70808 20547
rect 70728 20488 70808 20516
rect 70728 20476 70734 20488
rect 65797 20451 65855 20457
rect 65797 20417 65809 20451
rect 65843 20448 65855 20451
rect 66162 20448 66168 20460
rect 65843 20420 66024 20448
rect 65843 20417 65855 20420
rect 65797 20411 65855 20417
rect 1670 20340 1676 20392
rect 1728 20380 1734 20392
rect 65153 20383 65211 20389
rect 65153 20380 65165 20383
rect 1728 20352 65165 20380
rect 1728 20340 1734 20352
rect 65153 20349 65165 20352
rect 65199 20380 65211 20383
rect 65889 20383 65947 20389
rect 65889 20380 65901 20383
rect 65199 20352 65901 20380
rect 65199 20349 65211 20352
rect 65153 20343 65211 20349
rect 65889 20349 65901 20352
rect 65935 20349 65947 20383
rect 65889 20343 65947 20349
rect 64966 20272 64972 20324
rect 65024 20312 65030 20324
rect 65996 20312 66024 20420
rect 66088 20420 66168 20448
rect 66088 20389 66116 20420
rect 66162 20408 66168 20420
rect 66220 20448 66226 20460
rect 66220 20420 68784 20448
rect 66220 20408 66226 20420
rect 68756 20389 68784 20420
rect 68830 20408 68836 20460
rect 68888 20448 68894 20460
rect 69641 20451 69699 20457
rect 69641 20448 69653 20451
rect 68888 20420 69653 20448
rect 68888 20408 68894 20420
rect 69641 20417 69653 20420
rect 69687 20417 69699 20451
rect 69641 20411 69699 20417
rect 73709 20451 73767 20457
rect 73709 20417 73721 20451
rect 73755 20448 73767 20451
rect 74184 20448 74212 20547
rect 74626 20544 74632 20556
rect 74684 20544 74690 20596
rect 73755 20420 74212 20448
rect 74537 20451 74595 20457
rect 73755 20417 73767 20420
rect 73709 20411 73767 20417
rect 74537 20417 74549 20451
rect 74583 20448 74595 20451
rect 74902 20448 74908 20460
rect 74583 20420 74908 20448
rect 74583 20417 74595 20420
rect 74537 20411 74595 20417
rect 74902 20408 74908 20420
rect 74960 20408 74966 20460
rect 66073 20383 66131 20389
rect 66073 20349 66085 20383
rect 66119 20349 66131 20383
rect 66073 20343 66131 20349
rect 68741 20383 68799 20389
rect 68741 20349 68753 20383
rect 68787 20380 68799 20383
rect 69290 20380 69296 20392
rect 68787 20352 69296 20380
rect 68787 20349 68799 20352
rect 68741 20343 68799 20349
rect 69290 20340 69296 20352
rect 69348 20340 69354 20392
rect 69382 20340 69388 20392
rect 69440 20380 69446 20392
rect 69440 20352 69485 20380
rect 69440 20340 69446 20352
rect 70394 20340 70400 20392
rect 70452 20380 70458 20392
rect 74718 20380 74724 20392
rect 70452 20352 74724 20380
rect 70452 20340 70458 20352
rect 74718 20340 74724 20352
rect 74776 20340 74782 20392
rect 65024 20284 69152 20312
rect 65024 20272 65030 20284
rect 65426 20244 65432 20256
rect 65387 20216 65432 20244
rect 65426 20204 65432 20216
rect 65484 20204 65490 20256
rect 68189 20247 68247 20253
rect 68189 20213 68201 20247
rect 68235 20244 68247 20247
rect 69014 20244 69020 20256
rect 68235 20216 69020 20244
rect 68235 20213 68247 20216
rect 68189 20207 68247 20213
rect 69014 20204 69020 20216
rect 69072 20204 69078 20256
rect 69124 20244 69152 20284
rect 70026 20244 70032 20256
rect 69124 20216 70032 20244
rect 70026 20204 70032 20216
rect 70084 20204 70090 20256
rect 73525 20247 73583 20253
rect 73525 20213 73537 20247
rect 73571 20244 73583 20247
rect 73614 20244 73620 20256
rect 73571 20216 73620 20244
rect 73571 20213 73583 20216
rect 73525 20207 73583 20213
rect 73614 20204 73620 20216
rect 73672 20204 73678 20256
rect 1104 20154 118864 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 96374 20154
rect 96426 20102 96438 20154
rect 96490 20102 96502 20154
rect 96554 20102 96566 20154
rect 96618 20102 96630 20154
rect 96682 20102 118864 20154
rect 1104 20080 118864 20102
rect 64966 20040 64972 20052
rect 64927 20012 64972 20040
rect 64966 20000 64972 20012
rect 65024 20000 65030 20052
rect 68830 20040 68836 20052
rect 68791 20012 68836 20040
rect 68830 20000 68836 20012
rect 68888 20000 68894 20052
rect 74902 20040 74908 20052
rect 74863 20012 74908 20040
rect 74902 20000 74908 20012
rect 74960 20000 74966 20052
rect 68370 19904 68376 19916
rect 64846 19876 68376 19904
rect 63589 19839 63647 19845
rect 63589 19805 63601 19839
rect 63635 19836 63647 19839
rect 64846 19836 64874 19876
rect 68370 19864 68376 19876
rect 68428 19904 68434 19916
rect 69382 19904 69388 19916
rect 68428 19876 69388 19904
rect 68428 19864 68434 19876
rect 69382 19864 69388 19876
rect 69440 19904 69446 19916
rect 73525 19907 73583 19913
rect 73525 19904 73537 19907
rect 69440 19876 73537 19904
rect 69440 19864 69446 19876
rect 73525 19873 73537 19876
rect 73571 19873 73583 19907
rect 73525 19867 73583 19873
rect 69014 19836 69020 19848
rect 63635 19808 64874 19836
rect 68975 19808 69020 19836
rect 63635 19805 63647 19808
rect 63589 19799 63647 19805
rect 69014 19796 69020 19808
rect 69072 19796 69078 19848
rect 73614 19796 73620 19848
rect 73672 19836 73678 19848
rect 73781 19839 73839 19845
rect 73781 19836 73793 19839
rect 73672 19808 73793 19836
rect 73672 19796 73678 19808
rect 73781 19805 73793 19808
rect 73827 19805 73839 19839
rect 73781 19799 73839 19805
rect 63856 19771 63914 19777
rect 63856 19737 63868 19771
rect 63902 19768 63914 19771
rect 64230 19768 64236 19780
rect 63902 19740 64236 19768
rect 63902 19737 63914 19740
rect 63856 19731 63914 19737
rect 64230 19728 64236 19740
rect 64288 19728 64294 19780
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 64874 19700 64880 19712
rect 1728 19672 64880 19700
rect 1728 19660 1734 19672
rect 64874 19660 64880 19672
rect 64932 19660 64938 19712
rect 70854 19660 70860 19712
rect 70912 19700 70918 19712
rect 74920 19700 74948 20000
rect 70912 19672 74948 19700
rect 70912 19660 70918 19672
rect 1104 19610 118864 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 81014 19610
rect 81066 19558 81078 19610
rect 81130 19558 81142 19610
rect 81194 19558 81206 19610
rect 81258 19558 81270 19610
rect 81322 19558 111734 19610
rect 111786 19558 111798 19610
rect 111850 19558 111862 19610
rect 111914 19558 111926 19610
rect 111978 19558 111990 19610
rect 112042 19558 118864 19610
rect 1104 19536 118864 19558
rect 64230 19496 64236 19508
rect 64191 19468 64236 19496
rect 64230 19456 64236 19468
rect 64288 19456 64294 19508
rect 64874 19456 64880 19508
rect 64932 19496 64938 19508
rect 66073 19499 66131 19505
rect 66073 19496 66085 19499
rect 64932 19468 66085 19496
rect 64932 19456 64938 19468
rect 66073 19465 66085 19468
rect 66119 19465 66131 19499
rect 66073 19459 66131 19465
rect 66809 19499 66867 19505
rect 66809 19465 66821 19499
rect 66855 19465 66867 19499
rect 66809 19459 66867 19465
rect 69753 19499 69811 19505
rect 69753 19465 69765 19499
rect 69799 19465 69811 19499
rect 69753 19459 69811 19465
rect 71133 19499 71191 19505
rect 71133 19465 71145 19499
rect 71179 19496 71191 19499
rect 73890 19496 73896 19508
rect 71179 19468 73896 19496
rect 71179 19465 71191 19468
rect 71133 19459 71191 19465
rect 1670 19428 1676 19440
rect 1631 19400 1676 19428
rect 1670 19388 1676 19400
rect 1728 19388 1734 19440
rect 66824 19428 66852 19459
rect 68618 19431 68676 19437
rect 68618 19428 68630 19431
rect 65628 19400 66392 19428
rect 66824 19400 68630 19428
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 64417 19363 64475 19369
rect 64417 19329 64429 19363
rect 64463 19360 64475 19363
rect 65426 19360 65432 19372
rect 64463 19332 65432 19360
rect 64463 19329 64475 19332
rect 64417 19323 64475 19329
rect 65426 19320 65432 19332
rect 65484 19320 65490 19372
rect 65628 19233 65656 19400
rect 65981 19363 66039 19369
rect 65981 19329 65993 19363
rect 66027 19360 66039 19363
rect 66364 19360 66392 19400
rect 68618 19397 68630 19400
rect 68664 19397 68676 19431
rect 68618 19391 68676 19397
rect 69768 19428 69796 19459
rect 73890 19456 73896 19468
rect 73948 19456 73954 19508
rect 118050 19496 118056 19508
rect 118011 19468 118056 19496
rect 118050 19456 118056 19468
rect 118108 19456 118114 19508
rect 69768 19400 70992 19428
rect 66993 19363 67051 19369
rect 66993 19360 67005 19363
rect 66027 19332 66300 19360
rect 66364 19332 67005 19360
rect 66027 19329 66039 19332
rect 65981 19323 66039 19329
rect 66162 19292 66168 19304
rect 66123 19264 66168 19292
rect 66162 19252 66168 19264
rect 66220 19252 66226 19304
rect 66272 19292 66300 19332
rect 66993 19329 67005 19332
rect 67039 19329 67051 19363
rect 69768 19360 69796 19400
rect 66993 19323 67051 19329
rect 67100 19332 69796 19360
rect 67100 19292 67128 19332
rect 70026 19320 70032 19372
rect 70084 19360 70090 19372
rect 70673 19363 70731 19369
rect 70673 19360 70685 19363
rect 70084 19332 70685 19360
rect 70084 19320 70090 19332
rect 70673 19329 70685 19332
rect 70719 19329 70731 19363
rect 70854 19360 70860 19372
rect 70815 19332 70860 19360
rect 70673 19323 70731 19329
rect 70854 19320 70860 19332
rect 70912 19320 70918 19372
rect 70964 19369 70992 19400
rect 70949 19363 71007 19369
rect 70949 19329 70961 19363
rect 70995 19329 71007 19363
rect 117866 19360 117872 19372
rect 117827 19332 117872 19360
rect 70949 19323 71007 19329
rect 117866 19320 117872 19332
rect 117924 19320 117930 19372
rect 68370 19292 68376 19304
rect 66272 19264 67128 19292
rect 68331 19264 68376 19292
rect 68370 19252 68376 19264
rect 68428 19252 68434 19304
rect 65613 19227 65671 19233
rect 65613 19193 65625 19227
rect 65659 19193 65671 19227
rect 65613 19187 65671 19193
rect 70670 19156 70676 19168
rect 70631 19128 70676 19156
rect 70670 19116 70676 19128
rect 70728 19116 70734 19168
rect 1104 19066 118864 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 96374 19066
rect 96426 19014 96438 19066
rect 96490 19014 96502 19066
rect 96554 19014 96566 19066
rect 96618 19014 96630 19066
rect 96682 19014 118864 19066
rect 1104 18992 118864 19014
rect 57330 18680 57336 18692
rect 57291 18652 57336 18680
rect 57330 18640 57336 18652
rect 57388 18640 57394 18692
rect 57609 18615 57667 18621
rect 57609 18581 57621 18615
rect 57655 18612 57667 18615
rect 117866 18612 117872 18624
rect 57655 18584 117872 18612
rect 57655 18581 57667 18584
rect 57609 18575 57667 18581
rect 117866 18572 117872 18584
rect 117924 18572 117930 18624
rect 1104 18522 118864 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 81014 18522
rect 81066 18470 81078 18522
rect 81130 18470 81142 18522
rect 81194 18470 81206 18522
rect 81258 18470 81270 18522
rect 81322 18470 111734 18522
rect 111786 18470 111798 18522
rect 111850 18470 111862 18522
rect 111914 18470 111926 18522
rect 111978 18470 111990 18522
rect 112042 18470 118864 18522
rect 1104 18448 118864 18470
rect 117774 18272 117780 18284
rect 117735 18244 117780 18272
rect 117774 18232 117780 18244
rect 117832 18232 117838 18284
rect 117866 18068 117872 18080
rect 117827 18040 117872 18068
rect 117866 18028 117872 18040
rect 117924 18028 117930 18080
rect 1104 17978 118864 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 96374 17978
rect 96426 17926 96438 17978
rect 96490 17926 96502 17978
rect 96554 17926 96566 17978
rect 96618 17926 96630 17978
rect 96682 17926 118864 17978
rect 1104 17904 118864 17926
rect 1394 17660 1400 17672
rect 1355 17632 1400 17660
rect 1394 17620 1400 17632
rect 1452 17620 1458 17672
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 1762 17524 1768 17536
rect 1627 17496 1768 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 1762 17484 1768 17496
rect 1820 17484 1826 17536
rect 1104 17434 118864 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 81014 17434
rect 81066 17382 81078 17434
rect 81130 17382 81142 17434
rect 81194 17382 81206 17434
rect 81258 17382 81270 17434
rect 81322 17382 111734 17434
rect 111786 17382 111798 17434
rect 111850 17382 111862 17434
rect 111914 17382 111926 17434
rect 111978 17382 111990 17434
rect 112042 17382 118864 17434
rect 1104 17360 118864 17382
rect 1104 16890 118864 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 96374 16890
rect 96426 16838 96438 16890
rect 96490 16838 96502 16890
rect 96554 16838 96566 16890
rect 96618 16838 96630 16890
rect 96682 16838 118864 16890
rect 1104 16816 118864 16838
rect 1104 16346 118864 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 81014 16346
rect 81066 16294 81078 16346
rect 81130 16294 81142 16346
rect 81194 16294 81206 16346
rect 81258 16294 81270 16346
rect 81322 16294 111734 16346
rect 111786 16294 111798 16346
rect 111850 16294 111862 16346
rect 111914 16294 111926 16346
rect 111978 16294 111990 16346
rect 112042 16294 118864 16346
rect 1104 16272 118864 16294
rect 1104 15802 118864 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 96374 15802
rect 96426 15750 96438 15802
rect 96490 15750 96502 15802
rect 96554 15750 96566 15802
rect 96618 15750 96630 15802
rect 96682 15750 118864 15802
rect 1104 15728 118864 15750
rect 117774 15416 117780 15428
rect 117735 15388 117780 15416
rect 117774 15376 117780 15388
rect 117832 15376 117838 15428
rect 70486 15308 70492 15360
rect 70544 15348 70550 15360
rect 117869 15351 117927 15357
rect 117869 15348 117881 15351
rect 70544 15320 117881 15348
rect 70544 15308 70550 15320
rect 117869 15317 117881 15320
rect 117915 15317 117927 15351
rect 117869 15311 117927 15317
rect 1104 15258 118864 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 81014 15258
rect 81066 15206 81078 15258
rect 81130 15206 81142 15258
rect 81194 15206 81206 15258
rect 81258 15206 81270 15258
rect 81322 15206 111734 15258
rect 111786 15206 111798 15258
rect 111850 15206 111862 15258
rect 111914 15206 111926 15258
rect 111978 15206 111990 15258
rect 112042 15206 118864 15258
rect 1104 15184 118864 15206
rect 1104 14714 118864 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 96374 14714
rect 96426 14662 96438 14714
rect 96490 14662 96502 14714
rect 96554 14662 96566 14714
rect 96618 14662 96630 14714
rect 96682 14662 118864 14714
rect 1104 14640 118864 14662
rect 1302 14492 1308 14544
rect 1360 14532 1366 14544
rect 1486 14532 1492 14544
rect 1360 14504 1492 14532
rect 1360 14492 1366 14504
rect 1486 14492 1492 14504
rect 1544 14492 1550 14544
rect 1854 14328 1860 14340
rect 1815 14300 1860 14328
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 1104 14170 118864 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 81014 14170
rect 81066 14118 81078 14170
rect 81130 14118 81142 14170
rect 81194 14118 81206 14170
rect 81258 14118 81270 14170
rect 81322 14118 111734 14170
rect 111786 14118 111798 14170
rect 111850 14118 111862 14170
rect 111914 14118 111926 14170
rect 111978 14118 111990 14170
rect 112042 14118 118864 14170
rect 1104 14096 118864 14118
rect 1104 13626 118864 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 96374 13626
rect 96426 13574 96438 13626
rect 96490 13574 96502 13626
rect 96554 13574 96566 13626
rect 96618 13574 96630 13626
rect 96682 13574 118864 13626
rect 1104 13552 118864 13574
rect 1104 13082 118864 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 81014 13082
rect 81066 13030 81078 13082
rect 81130 13030 81142 13082
rect 81194 13030 81206 13082
rect 81258 13030 81270 13082
rect 81322 13030 111734 13082
rect 111786 13030 111798 13082
rect 111850 13030 111862 13082
rect 111914 13030 111926 13082
rect 111978 13030 111990 13082
rect 112042 13030 118864 13082
rect 1104 13008 118864 13030
rect 1104 12538 118864 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 96374 12538
rect 96426 12486 96438 12538
rect 96490 12486 96502 12538
rect 96554 12486 96566 12538
rect 96618 12486 96630 12538
rect 96682 12486 118864 12538
rect 1104 12464 118864 12486
rect 117222 12152 117228 12164
rect 117183 12124 117228 12152
rect 117222 12112 117228 12124
rect 117280 12112 117286 12164
rect 117961 12155 118019 12161
rect 117961 12121 117973 12155
rect 118007 12121 118019 12155
rect 117961 12115 118019 12121
rect 39666 12044 39672 12096
rect 39724 12084 39730 12096
rect 117976 12084 118004 12115
rect 39724 12056 118004 12084
rect 39724 12044 39730 12056
rect 1104 11994 118864 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 81014 11994
rect 81066 11942 81078 11994
rect 81130 11942 81142 11994
rect 81194 11942 81206 11994
rect 81258 11942 81270 11994
rect 81322 11942 111734 11994
rect 111786 11942 111798 11994
rect 111850 11942 111862 11994
rect 111914 11942 111926 11994
rect 111978 11942 111990 11994
rect 112042 11942 118864 11994
rect 1104 11920 118864 11942
rect 1104 11450 118864 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 96374 11450
rect 96426 11398 96438 11450
rect 96490 11398 96502 11450
rect 96554 11398 96566 11450
rect 96618 11398 96630 11450
rect 96682 11398 118864 11450
rect 1104 11376 118864 11398
rect 1854 11064 1860 11076
rect 1815 11036 1860 11064
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2041 11067 2099 11073
rect 2041 11033 2053 11067
rect 2087 11064 2099 11067
rect 7558 11064 7564 11076
rect 2087 11036 7564 11064
rect 2087 11033 2099 11036
rect 2041 11027 2099 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 1104 10906 118864 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 81014 10906
rect 81066 10854 81078 10906
rect 81130 10854 81142 10906
rect 81194 10854 81206 10906
rect 81258 10854 81270 10906
rect 81322 10854 111734 10906
rect 111786 10854 111798 10906
rect 111850 10854 111862 10906
rect 111914 10854 111926 10906
rect 111978 10854 111990 10906
rect 112042 10854 118864 10906
rect 1104 10832 118864 10854
rect 1854 10684 1860 10736
rect 1912 10724 1918 10736
rect 2038 10724 2044 10736
rect 1912 10696 2044 10724
rect 1912 10684 1918 10696
rect 2038 10684 2044 10696
rect 2096 10684 2102 10736
rect 1104 10362 118864 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 96374 10362
rect 96426 10310 96438 10362
rect 96490 10310 96502 10362
rect 96554 10310 96566 10362
rect 96618 10310 96630 10362
rect 96682 10310 118864 10362
rect 1104 10288 118864 10310
rect 1104 9818 118864 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 81014 9818
rect 81066 9766 81078 9818
rect 81130 9766 81142 9818
rect 81194 9766 81206 9818
rect 81258 9766 81270 9818
rect 81322 9766 111734 9818
rect 111786 9766 111798 9818
rect 111850 9766 111862 9818
rect 111914 9766 111926 9818
rect 111978 9766 111990 9818
rect 112042 9766 118864 9818
rect 1104 9744 118864 9766
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9568 1455 9571
rect 22094 9568 22100 9580
rect 1443 9540 22100 9568
rect 1443 9537 1455 9540
rect 1397 9531 1455 9537
rect 22094 9528 22100 9540
rect 22152 9528 22158 9580
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1104 9274 118864 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 96374 9274
rect 96426 9222 96438 9274
rect 96490 9222 96502 9274
rect 96554 9222 96566 9274
rect 96618 9222 96630 9274
rect 96682 9222 118864 9274
rect 1104 9200 118864 9222
rect 1104 8730 118864 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 81014 8730
rect 81066 8678 81078 8730
rect 81130 8678 81142 8730
rect 81194 8678 81206 8730
rect 81258 8678 81270 8730
rect 81322 8678 111734 8730
rect 111786 8678 111798 8730
rect 111850 8678 111862 8730
rect 111914 8678 111926 8730
rect 111978 8678 111990 8730
rect 112042 8678 118864 8730
rect 1104 8656 118864 8678
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8480 21879 8483
rect 22370 8480 22376 8492
rect 21867 8452 22376 8480
rect 21867 8449 21879 8452
rect 21821 8443 21879 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22094 8412 22100 8424
rect 22055 8384 22100 8412
rect 22094 8372 22100 8384
rect 22152 8372 22158 8424
rect 1104 8186 118864 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 96374 8186
rect 96426 8134 96438 8186
rect 96490 8134 96502 8186
rect 96554 8134 96566 8186
rect 96618 8134 96630 8186
rect 96682 8134 118864 8186
rect 1104 8112 118864 8134
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 10318 7732 10324 7744
rect 1443 7704 10324 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 1104 7642 118864 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 81014 7642
rect 81066 7590 81078 7642
rect 81130 7590 81142 7642
rect 81194 7590 81206 7642
rect 81258 7590 81270 7642
rect 81322 7590 111734 7642
rect 111786 7590 111798 7642
rect 111850 7590 111862 7642
rect 111914 7590 111926 7642
rect 111978 7590 111990 7642
rect 112042 7590 118864 7642
rect 1104 7568 118864 7590
rect 1104 7098 118864 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 118864 7098
rect 1104 7024 118864 7046
rect 117958 6712 117964 6724
rect 117919 6684 117964 6712
rect 117958 6672 117964 6684
rect 118016 6672 118022 6724
rect 114462 6604 114468 6656
rect 114520 6644 114526 6656
rect 118053 6647 118111 6653
rect 118053 6644 118065 6647
rect 114520 6616 118065 6644
rect 114520 6604 114526 6616
rect 118053 6613 118065 6616
rect 118099 6613 118111 6647
rect 118053 6607 118111 6613
rect 1104 6554 118864 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 81014 6554
rect 81066 6502 81078 6554
rect 81130 6502 81142 6554
rect 81194 6502 81206 6554
rect 81258 6502 81270 6554
rect 81322 6502 111734 6554
rect 111786 6502 111798 6554
rect 111850 6502 111862 6554
rect 111914 6502 111926 6554
rect 111978 6502 111990 6554
rect 112042 6502 118864 6554
rect 1104 6480 118864 6502
rect 76653 6443 76711 6449
rect 76653 6409 76665 6443
rect 76699 6409 76711 6443
rect 77110 6440 77116 6452
rect 77071 6412 77116 6440
rect 76653 6403 76711 6409
rect 76009 6307 76067 6313
rect 76009 6273 76021 6307
rect 76055 6304 76067 6307
rect 76668 6304 76696 6403
rect 77110 6400 77116 6412
rect 77168 6400 77174 6452
rect 76055 6276 76696 6304
rect 76055 6273 76067 6276
rect 76009 6267 76067 6273
rect 76926 6264 76932 6316
rect 76984 6304 76990 6316
rect 77021 6307 77079 6313
rect 77021 6304 77033 6307
rect 76984 6276 77033 6304
rect 76984 6264 76990 6276
rect 77021 6273 77033 6276
rect 77067 6273 77079 6307
rect 77021 6267 77079 6273
rect 77202 6236 77208 6248
rect 77163 6208 77208 6236
rect 77202 6196 77208 6208
rect 77260 6196 77266 6248
rect 75825 6103 75883 6109
rect 75825 6069 75837 6103
rect 75871 6100 75883 6103
rect 76006 6100 76012 6112
rect 75871 6072 76012 6100
rect 75871 6069 75883 6072
rect 75825 6063 75883 6069
rect 76006 6060 76012 6072
rect 76064 6060 76070 6112
rect 1104 6010 118864 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 118864 6010
rect 1104 5936 118864 5958
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 17218 5692 17224 5704
rect 17179 5664 17224 5692
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 75914 5692 75920 5704
rect 75875 5664 75920 5692
rect 75914 5652 75920 5664
rect 75972 5652 75978 5704
rect 76006 5652 76012 5704
rect 76064 5692 76070 5704
rect 76173 5695 76231 5701
rect 76173 5692 76185 5695
rect 76064 5664 76185 5692
rect 76064 5652 76070 5664
rect 76173 5661 76185 5664
rect 76219 5661 76231 5695
rect 76173 5655 76231 5661
rect 9858 5556 9864 5568
rect 9819 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 17037 5559 17095 5565
rect 17037 5525 17049 5559
rect 17083 5556 17095 5559
rect 17126 5556 17132 5568
rect 17083 5528 17132 5556
rect 17083 5525 17095 5528
rect 17037 5519 17095 5525
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 76926 5516 76932 5568
rect 76984 5556 76990 5568
rect 77297 5559 77355 5565
rect 77297 5556 77309 5559
rect 76984 5528 77309 5556
rect 76984 5516 76990 5528
rect 77297 5525 77309 5528
rect 77343 5525 77355 5559
rect 77297 5519 77355 5525
rect 1104 5466 118864 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 81014 5466
rect 81066 5414 81078 5466
rect 81130 5414 81142 5466
rect 81194 5414 81206 5466
rect 81258 5414 81270 5466
rect 81322 5414 111734 5466
rect 111786 5414 111798 5466
rect 111850 5414 111862 5466
rect 111914 5414 111926 5466
rect 111978 5414 111990 5466
rect 112042 5414 118864 5466
rect 1104 5392 118864 5414
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10042 5352 10048 5364
rect 9907 5324 10048 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 10318 5352 10324 5364
rect 10279 5324 10324 5352
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17218 5352 17224 5364
rect 17175 5324 17224 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 27893 5355 27951 5361
rect 27893 5352 27905 5355
rect 20864 5324 27905 5352
rect 20864 5312 20870 5324
rect 27893 5321 27905 5324
rect 27939 5352 27951 5355
rect 28721 5355 28779 5361
rect 28721 5352 28733 5355
rect 27939 5324 28733 5352
rect 27939 5321 27951 5324
rect 27893 5315 27951 5321
rect 28721 5321 28733 5324
rect 28767 5321 28779 5355
rect 28721 5315 28779 5321
rect 39209 5355 39267 5361
rect 39209 5321 39221 5355
rect 39255 5321 39267 5355
rect 39666 5352 39672 5364
rect 39627 5324 39672 5352
rect 39209 5315 39267 5321
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 17589 5287 17647 5293
rect 17589 5284 17601 5287
rect 7616 5256 17601 5284
rect 7616 5244 7622 5256
rect 17589 5253 17601 5256
rect 17635 5253 17647 5287
rect 17589 5247 17647 5253
rect 20732 5256 22508 5284
rect 10226 5216 10232 5228
rect 10187 5188 10232 5216
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 18414 5216 18420 5228
rect 17543 5188 18420 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 18414 5176 18420 5188
rect 18472 5176 18478 5228
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 10551 5120 17785 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 17773 5117 17785 5120
rect 17819 5148 17831 5151
rect 20732 5148 20760 5256
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 22186 5216 22192 5228
rect 21315 5188 21864 5216
rect 22147 5188 22192 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 17819 5120 20760 5148
rect 17819 5117 17831 5120
rect 17773 5111 17831 5117
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 21836 5089 21864 5188
rect 22186 5176 22192 5188
rect 22244 5176 22250 5228
rect 22480 5157 22508 5256
rect 28626 5216 28632 5228
rect 28587 5188 28632 5216
rect 28626 5176 28632 5188
rect 28684 5176 28690 5228
rect 38749 5219 38807 5225
rect 38749 5185 38761 5219
rect 38795 5216 38807 5219
rect 39224 5216 39252 5315
rect 39666 5312 39672 5324
rect 39724 5312 39730 5364
rect 39850 5312 39856 5364
rect 39908 5352 39914 5364
rect 49878 5352 49884 5364
rect 39908 5324 49884 5352
rect 39908 5312 39914 5324
rect 49878 5312 49884 5324
rect 49936 5312 49942 5364
rect 49970 5312 49976 5364
rect 50028 5352 50034 5364
rect 50062 5352 50068 5364
rect 50028 5324 50068 5352
rect 50028 5312 50034 5324
rect 50062 5312 50068 5324
rect 50120 5352 50126 5364
rect 50890 5352 50896 5364
rect 50120 5324 50384 5352
rect 50851 5324 50896 5352
rect 50120 5312 50126 5324
rect 50356 5284 50384 5324
rect 50890 5312 50896 5324
rect 50948 5312 50954 5364
rect 63957 5355 64015 5361
rect 63957 5321 63969 5355
rect 64003 5321 64015 5355
rect 64414 5352 64420 5364
rect 64375 5324 64420 5352
rect 63957 5315 64015 5321
rect 50801 5287 50859 5293
rect 50801 5284 50813 5287
rect 48286 5256 50016 5284
rect 50356 5256 50813 5284
rect 39574 5216 39580 5228
rect 38795 5188 39252 5216
rect 39535 5188 39580 5216
rect 38795 5185 38807 5188
rect 38749 5179 38807 5185
rect 39574 5176 39580 5188
rect 39632 5176 39638 5228
rect 48286 5216 48314 5256
rect 39684 5188 48314 5216
rect 48860 5219 48918 5225
rect 22281 5151 22339 5157
rect 22281 5117 22293 5151
rect 22327 5117 22339 5151
rect 22281 5111 22339 5117
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 28905 5151 28963 5157
rect 22511 5120 26234 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 21821 5083 21879 5089
rect 2004 5052 21772 5080
rect 2004 5040 2010 5052
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 20806 5012 20812 5024
rect 1820 4984 20812 5012
rect 1820 4972 1826 4984
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 21085 5015 21143 5021
rect 21085 4981 21097 5015
rect 21131 5012 21143 5015
rect 21358 5012 21364 5024
rect 21131 4984 21364 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 21744 5012 21772 5052
rect 21821 5049 21833 5083
rect 21867 5049 21879 5083
rect 21821 5043 21879 5049
rect 22296 5080 22324 5111
rect 22833 5083 22891 5089
rect 22833 5080 22845 5083
rect 22296 5052 22845 5080
rect 22296 5012 22324 5052
rect 22833 5049 22845 5052
rect 22879 5049 22891 5083
rect 26206 5080 26234 5120
rect 28905 5117 28917 5151
rect 28951 5148 28963 5151
rect 39684 5148 39712 5188
rect 48860 5185 48872 5219
rect 48906 5216 48918 5219
rect 49326 5216 49332 5228
rect 48906 5188 49332 5216
rect 48906 5185 48918 5188
rect 48860 5179 48918 5185
rect 49326 5176 49332 5188
rect 49384 5176 49390 5228
rect 49988 5216 50016 5256
rect 50801 5253 50813 5256
rect 50847 5253 50859 5287
rect 50801 5247 50859 5253
rect 49988 5188 53328 5216
rect 39850 5148 39856 5160
rect 28951 5120 39712 5148
rect 39811 5120 39856 5148
rect 28951 5117 28963 5120
rect 28905 5111 28963 5117
rect 39850 5108 39856 5120
rect 39908 5108 39914 5160
rect 48590 5148 48596 5160
rect 48551 5120 48596 5148
rect 48590 5108 48596 5120
rect 48648 5108 48654 5160
rect 49878 5108 49884 5160
rect 49936 5148 49942 5160
rect 50982 5148 50988 5160
rect 49936 5120 50988 5148
rect 49936 5108 49942 5120
rect 50982 5108 50988 5120
rect 51040 5108 51046 5160
rect 53300 5148 53328 5188
rect 53558 5176 53564 5228
rect 53616 5216 53622 5228
rect 63221 5219 63279 5225
rect 53616 5188 53661 5216
rect 53616 5176 53622 5188
rect 63221 5185 63233 5219
rect 63267 5216 63279 5219
rect 63972 5216 64000 5315
rect 64414 5312 64420 5324
rect 64472 5312 64478 5364
rect 70029 5355 70087 5361
rect 70029 5321 70041 5355
rect 70075 5321 70087 5355
rect 70486 5352 70492 5364
rect 70447 5324 70492 5352
rect 70029 5315 70087 5321
rect 63267 5188 64000 5216
rect 63267 5185 63279 5188
rect 63221 5179 63279 5185
rect 64046 5176 64052 5228
rect 64104 5216 64110 5228
rect 64325 5219 64383 5225
rect 64325 5216 64337 5219
rect 64104 5188 64337 5216
rect 64104 5176 64110 5188
rect 64325 5185 64337 5188
rect 64371 5185 64383 5219
rect 64325 5179 64383 5185
rect 68741 5219 68799 5225
rect 68741 5185 68753 5219
rect 68787 5216 68799 5219
rect 70044 5216 70072 5315
rect 70486 5312 70492 5324
rect 70544 5312 70550 5364
rect 75825 5355 75883 5361
rect 75825 5352 75837 5355
rect 73632 5324 75837 5352
rect 68787 5188 70072 5216
rect 68787 5185 68799 5188
rect 68741 5179 68799 5185
rect 70118 5176 70124 5228
rect 70176 5216 70182 5228
rect 73632 5225 73660 5324
rect 75825 5321 75837 5324
rect 75871 5321 75883 5355
rect 92014 5352 92020 5364
rect 91975 5324 92020 5352
rect 75825 5315 75883 5321
rect 92014 5312 92020 5324
rect 92072 5312 92078 5364
rect 97626 5312 97632 5364
rect 97684 5352 97690 5364
rect 100665 5355 100723 5361
rect 100665 5352 100677 5355
rect 97684 5324 100677 5352
rect 97684 5312 97690 5324
rect 100665 5321 100677 5324
rect 100711 5352 100723 5355
rect 103790 5352 103796 5364
rect 100711 5324 103796 5352
rect 100711 5321 100723 5324
rect 100665 5315 100723 5321
rect 103790 5312 103796 5324
rect 103848 5312 103854 5364
rect 106752 5324 109034 5352
rect 74442 5244 74448 5296
rect 74500 5284 74506 5296
rect 76193 5287 76251 5293
rect 76193 5284 76205 5287
rect 74500 5256 76205 5284
rect 74500 5244 74506 5256
rect 76193 5253 76205 5256
rect 76239 5253 76251 5287
rect 76193 5247 76251 5253
rect 76285 5287 76343 5293
rect 76285 5253 76297 5287
rect 76331 5284 76343 5287
rect 106752 5284 106780 5324
rect 76331 5256 102732 5284
rect 76331 5253 76343 5256
rect 76285 5247 76343 5253
rect 70397 5219 70455 5225
rect 70397 5216 70409 5219
rect 70176 5188 70409 5216
rect 70176 5176 70182 5188
rect 70397 5185 70409 5188
rect 70443 5185 70455 5219
rect 70397 5179 70455 5185
rect 73617 5219 73675 5225
rect 73617 5185 73629 5219
rect 73663 5185 73675 5219
rect 73617 5179 73675 5185
rect 75549 5219 75607 5225
rect 75549 5185 75561 5219
rect 75595 5216 75607 5219
rect 76300 5216 76328 5247
rect 91922 5216 91928 5228
rect 75595 5188 76328 5216
rect 91883 5188 91928 5216
rect 75595 5185 75607 5188
rect 75549 5179 75607 5185
rect 91922 5176 91928 5188
rect 91980 5176 91986 5228
rect 96798 5216 96804 5228
rect 96724 5188 96804 5216
rect 53745 5151 53803 5157
rect 53745 5148 53757 5151
rect 53300 5120 53757 5148
rect 53745 5117 53757 5120
rect 53791 5148 53803 5151
rect 64509 5151 64567 5157
rect 64509 5148 64521 5151
rect 53791 5120 64521 5148
rect 53791 5117 53803 5120
rect 53745 5111 53803 5117
rect 64509 5117 64521 5120
rect 64555 5148 64567 5151
rect 70581 5151 70639 5157
rect 70581 5148 70593 5151
rect 64555 5120 70593 5148
rect 64555 5117 64567 5120
rect 64509 5111 64567 5117
rect 70581 5117 70593 5120
rect 70627 5148 70639 5151
rect 76377 5151 76435 5157
rect 70627 5120 74534 5148
rect 70627 5117 70639 5120
rect 70581 5111 70639 5117
rect 39868 5080 39896 5108
rect 61654 5080 61660 5092
rect 26206 5052 39896 5080
rect 49528 5052 61660 5080
rect 22833 5043 22891 5049
rect 21744 4984 22324 5012
rect 28261 5015 28319 5021
rect 28261 4981 28273 5015
rect 28307 5012 28319 5015
rect 29730 5012 29736 5024
rect 28307 4984 29736 5012
rect 28307 4981 28319 4984
rect 28261 4975 28319 4981
rect 29730 4972 29736 4984
rect 29788 4972 29794 5024
rect 38565 5015 38623 5021
rect 38565 4981 38577 5015
rect 38611 5012 38623 5015
rect 38654 5012 38660 5024
rect 38611 4984 38660 5012
rect 38611 4981 38623 4984
rect 38565 4975 38623 4981
rect 38654 4972 38660 4984
rect 38712 4972 38718 5024
rect 48590 4972 48596 5024
rect 48648 5012 48654 5024
rect 49528 5012 49556 5052
rect 61654 5040 61660 5052
rect 61712 5040 61718 5092
rect 74506 5080 74534 5120
rect 76377 5117 76389 5151
rect 76423 5148 76435 5151
rect 77202 5148 77208 5160
rect 76423 5120 77208 5148
rect 76423 5117 76435 5120
rect 76377 5111 76435 5117
rect 76392 5080 76420 5111
rect 77202 5108 77208 5120
rect 77260 5108 77266 5160
rect 92109 5151 92167 5157
rect 92109 5117 92121 5151
rect 92155 5117 92167 5151
rect 92109 5111 92167 5117
rect 74506 5052 76420 5080
rect 77294 5040 77300 5092
rect 77352 5080 77358 5092
rect 92124 5080 92152 5111
rect 94038 5108 94044 5160
rect 94096 5148 94102 5160
rect 96724 5157 96752 5188
rect 96798 5176 96804 5188
rect 96856 5176 96862 5228
rect 96982 5225 96988 5228
rect 96976 5179 96988 5225
rect 97040 5216 97046 5228
rect 100754 5216 100760 5228
rect 97040 5188 97076 5216
rect 100715 5188 100760 5216
rect 96982 5176 96988 5179
rect 97040 5176 97046 5188
rect 100754 5176 100760 5188
rect 100812 5176 100818 5228
rect 102577 5219 102635 5225
rect 102577 5216 102589 5219
rect 101508 5188 102589 5216
rect 96709 5151 96767 5157
rect 96709 5148 96721 5151
rect 94096 5120 96721 5148
rect 94096 5108 94102 5120
rect 96709 5117 96721 5120
rect 96755 5117 96767 5151
rect 100294 5148 100300 5160
rect 100255 5120 100300 5148
rect 96709 5111 96767 5117
rect 100294 5108 100300 5120
rect 100352 5108 100358 5160
rect 100481 5151 100539 5157
rect 100481 5117 100493 5151
rect 100527 5148 100539 5151
rect 101508 5148 101536 5188
rect 102577 5185 102589 5188
rect 102623 5185 102635 5219
rect 102704 5216 102732 5256
rect 103900 5256 106780 5284
rect 109006 5284 109034 5324
rect 117774 5284 117780 5296
rect 109006 5256 117780 5284
rect 103900 5216 103928 5256
rect 117774 5244 117780 5256
rect 117832 5244 117838 5296
rect 102704 5188 103928 5216
rect 102577 5179 102635 5185
rect 104526 5176 104532 5228
rect 104584 5216 104590 5228
rect 106717 5219 106775 5225
rect 106717 5216 106729 5219
rect 104584 5188 106729 5216
rect 104584 5176 104590 5188
rect 106717 5185 106729 5188
rect 106763 5185 106775 5219
rect 117869 5219 117927 5225
rect 106717 5179 106775 5185
rect 109006 5188 113174 5216
rect 102318 5148 102324 5160
rect 100527 5120 101536 5148
rect 102279 5120 102324 5148
rect 100527 5117 100539 5120
rect 100481 5111 100539 5117
rect 102318 5108 102324 5120
rect 102376 5108 102382 5160
rect 106458 5148 106464 5160
rect 106419 5120 106464 5148
rect 106458 5108 106464 5120
rect 106516 5108 106522 5160
rect 96614 5080 96620 5092
rect 77352 5052 96620 5080
rect 77352 5040 77358 5052
rect 96614 5040 96620 5052
rect 96672 5040 96678 5092
rect 109006 5080 109034 5188
rect 107396 5052 109034 5080
rect 113146 5080 113174 5188
rect 117869 5185 117881 5219
rect 117915 5185 117927 5219
rect 117869 5179 117927 5185
rect 114462 5080 114468 5092
rect 113146 5052 114468 5080
rect 48648 4984 49556 5012
rect 48648 4972 48654 4984
rect 50062 4972 50068 5024
rect 50120 5012 50126 5024
rect 50433 5015 50491 5021
rect 50433 5012 50445 5015
rect 50120 4984 50445 5012
rect 50120 4972 50126 4984
rect 50433 4981 50445 4984
rect 50479 4981 50491 5015
rect 63034 5012 63040 5024
rect 62995 4984 63040 5012
rect 50433 4975 50491 4981
rect 63034 4972 63040 4984
rect 63092 4972 63098 5024
rect 68554 5012 68560 5024
rect 68515 4984 68560 5012
rect 68554 4972 68560 4984
rect 68612 4972 68618 5024
rect 73430 5012 73436 5024
rect 73391 4984 73436 5012
rect 73430 4972 73436 4984
rect 73488 4972 73494 5024
rect 91094 4972 91100 5024
rect 91152 5012 91158 5024
rect 91557 5015 91615 5021
rect 91557 5012 91569 5015
rect 91152 4984 91569 5012
rect 91152 4972 91158 4984
rect 91557 4981 91569 4984
rect 91603 4981 91615 5015
rect 91557 4975 91615 4981
rect 93946 4972 93952 5024
rect 94004 5012 94010 5024
rect 98089 5015 98147 5021
rect 98089 5012 98101 5015
rect 94004 4984 98101 5012
rect 94004 4972 94010 4984
rect 98089 4981 98101 4984
rect 98135 5012 98147 5015
rect 100202 5012 100208 5024
rect 98135 4984 100208 5012
rect 98135 4981 98147 4984
rect 98089 4975 98147 4981
rect 100202 4972 100208 4984
rect 100260 4972 100266 5024
rect 100938 4972 100944 5024
rect 100996 5012 101002 5024
rect 103701 5015 103759 5021
rect 103701 5012 103713 5015
rect 100996 4984 103713 5012
rect 100996 4972 101002 4984
rect 103701 4981 103713 4984
rect 103747 4981 103759 5015
rect 103701 4975 103759 4981
rect 103790 4972 103796 5024
rect 103848 5012 103854 5024
rect 107396 5012 107424 5052
rect 114462 5040 114468 5052
rect 114520 5040 114526 5092
rect 107838 5012 107844 5024
rect 103848 4984 107424 5012
rect 107799 4984 107844 5012
rect 103848 4972 103854 4984
rect 107838 4972 107844 4984
rect 107896 5012 107902 5024
rect 117884 5012 117912 5179
rect 118050 5012 118056 5024
rect 107896 4984 117912 5012
rect 118011 4984 118056 5012
rect 107896 4972 107902 4984
rect 118050 4972 118056 4984
rect 118108 4972 118114 5024
rect 1104 4922 118864 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 118864 4922
rect 1104 4848 118864 4870
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 22186 4768 22192 4820
rect 22244 4808 22250 4820
rect 22649 4811 22707 4817
rect 22649 4808 22661 4811
rect 22244 4780 22661 4808
rect 22244 4768 22250 4780
rect 22649 4777 22661 4780
rect 22695 4808 22707 4811
rect 22738 4808 22744 4820
rect 22695 4780 22744 4808
rect 22695 4777 22707 4780
rect 22649 4771 22707 4777
rect 22738 4768 22744 4780
rect 22796 4768 22802 4820
rect 38562 4808 38568 4820
rect 27540 4780 38568 4808
rect 27540 4681 27568 4780
rect 38562 4768 38568 4780
rect 38620 4808 38626 4820
rect 48590 4808 48596 4820
rect 38620 4780 48596 4808
rect 38620 4768 38626 4780
rect 48590 4768 48596 4780
rect 48648 4768 48654 4820
rect 49326 4808 49332 4820
rect 49287 4780 49332 4808
rect 49326 4768 49332 4780
rect 49384 4768 49390 4820
rect 63037 4811 63095 4817
rect 63037 4777 63049 4811
rect 63083 4808 63095 4811
rect 63126 4808 63132 4820
rect 63083 4780 63132 4808
rect 63083 4777 63095 4780
rect 63037 4771 63095 4777
rect 63126 4768 63132 4780
rect 63184 4808 63190 4820
rect 64046 4808 64052 4820
rect 63184 4780 64052 4808
rect 63184 4768 63190 4780
rect 64046 4768 64052 4780
rect 64104 4768 64110 4820
rect 69198 4808 69204 4820
rect 69111 4780 69204 4808
rect 69198 4768 69204 4780
rect 69256 4808 69262 4820
rect 70118 4808 70124 4820
rect 69256 4780 70124 4808
rect 69256 4768 69262 4780
rect 70118 4768 70124 4780
rect 70176 4768 70182 4820
rect 76926 4808 76932 4820
rect 76887 4780 76932 4808
rect 76926 4768 76932 4780
rect 76984 4768 76990 4820
rect 90821 4811 90879 4817
rect 90821 4777 90833 4811
rect 90867 4808 90879 4811
rect 91922 4808 91928 4820
rect 90867 4780 91928 4808
rect 90867 4777 90879 4780
rect 90821 4771 90879 4777
rect 91922 4768 91928 4780
rect 91980 4768 91986 4820
rect 96982 4768 96988 4820
rect 97040 4808 97046 4820
rect 97169 4811 97227 4817
rect 97169 4808 97181 4811
rect 97040 4780 97181 4808
rect 97040 4768 97046 4780
rect 97169 4777 97181 4780
rect 97215 4777 97227 4811
rect 97169 4771 97227 4777
rect 100205 4811 100263 4817
rect 100205 4777 100217 4811
rect 100251 4808 100263 4811
rect 100754 4808 100760 4820
rect 100251 4780 100760 4808
rect 100251 4777 100263 4780
rect 100205 4771 100263 4777
rect 100754 4768 100760 4780
rect 100812 4768 100818 4820
rect 104526 4808 104532 4820
rect 104487 4780 104532 4808
rect 104526 4768 104532 4780
rect 104584 4768 104590 4820
rect 75914 4700 75920 4752
rect 75972 4740 75978 4752
rect 86218 4740 86224 4752
rect 75972 4712 86224 4740
rect 75972 4700 75978 4712
rect 86218 4700 86224 4712
rect 86276 4700 86282 4752
rect 100294 4740 100300 4752
rect 97460 4712 100300 4740
rect 27525 4675 27583 4681
rect 27525 4641 27537 4675
rect 27571 4641 27583 4675
rect 27525 4635 27583 4641
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 2464 4576 9597 4604
rect 2464 4564 2470 4576
rect 9585 4573 9597 4576
rect 9631 4604 9643 4607
rect 17037 4607 17095 4613
rect 17037 4604 17049 4607
rect 9631 4576 17049 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 17037 4573 17049 4576
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 9858 4545 9864 4548
rect 9852 4536 9864 4545
rect 9819 4508 9864 4536
rect 9852 4499 9864 4508
rect 9858 4496 9864 4499
rect 9916 4496 9922 4548
rect 17052 4536 17080 4567
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 17293 4607 17351 4613
rect 17293 4604 17305 4607
rect 17184 4576 17305 4604
rect 17184 4564 17190 4576
rect 17293 4573 17305 4576
rect 17339 4573 17351 4607
rect 17293 4567 17351 4573
rect 21269 4607 21327 4613
rect 21269 4573 21281 4607
rect 21315 4573 21327 4607
rect 21269 4567 21327 4573
rect 21284 4536 21312 4567
rect 21358 4564 21364 4616
rect 21416 4604 21422 4616
rect 21525 4607 21583 4613
rect 21525 4604 21537 4607
rect 21416 4576 21537 4604
rect 21416 4564 21422 4576
rect 21525 4573 21537 4576
rect 21571 4573 21583 4607
rect 21525 4567 21583 4573
rect 27540 4536 27568 4635
rect 49970 4632 49976 4684
rect 50028 4672 50034 4684
rect 50157 4675 50215 4681
rect 50157 4672 50169 4675
rect 50028 4644 50169 4672
rect 50028 4632 50034 4644
rect 50157 4641 50169 4644
rect 50203 4641 50215 4675
rect 50157 4635 50215 4641
rect 50982 4632 50988 4684
rect 51040 4672 51046 4684
rect 52733 4675 52791 4681
rect 52733 4672 52745 4675
rect 51040 4644 52745 4672
rect 51040 4632 51046 4644
rect 52733 4641 52745 4644
rect 52779 4641 52791 4675
rect 61654 4672 61660 4684
rect 61615 4644 61660 4672
rect 52733 4635 52791 4641
rect 61654 4632 61660 4644
rect 61712 4632 61718 4684
rect 73982 4632 73988 4684
rect 74040 4672 74046 4684
rect 76745 4675 76803 4681
rect 76745 4672 76757 4675
rect 74040 4644 76757 4672
rect 74040 4632 74046 4644
rect 76745 4641 76757 4644
rect 76791 4641 76803 4675
rect 86236 4672 86264 4700
rect 89441 4675 89499 4681
rect 89441 4672 89453 4675
rect 86236 4644 89453 4672
rect 76745 4635 76803 4641
rect 89441 4641 89453 4644
rect 89487 4641 89499 4675
rect 89441 4635 89499 4641
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 49513 4607 49571 4613
rect 49513 4573 49525 4607
rect 49559 4604 49571 4607
rect 50062 4604 50068 4616
rect 49559 4576 50068 4604
rect 49559 4573 49571 4576
rect 49513 4567 49571 4573
rect 50062 4564 50068 4576
rect 50120 4564 50126 4616
rect 50341 4607 50399 4613
rect 50341 4573 50353 4607
rect 50387 4604 50399 4607
rect 50614 4604 50620 4616
rect 50387 4576 50620 4604
rect 50387 4573 50399 4576
rect 50341 4567 50399 4573
rect 50614 4564 50620 4576
rect 50672 4564 50678 4616
rect 52549 4607 52607 4613
rect 52549 4573 52561 4607
rect 52595 4604 52607 4607
rect 53558 4604 53564 4616
rect 52595 4576 53564 4604
rect 52595 4573 52607 4576
rect 52549 4567 52607 4573
rect 53558 4564 53564 4576
rect 53616 4564 53622 4616
rect 17052 4508 27568 4536
rect 27792 4539 27850 4545
rect 27792 4505 27804 4539
rect 27838 4536 27850 4539
rect 61672 4536 61700 4632
rect 61924 4607 61982 4613
rect 61924 4573 61936 4607
rect 61970 4604 61982 4607
rect 63034 4604 63040 4616
rect 61970 4576 63040 4604
rect 61970 4573 61982 4576
rect 61924 4567 61982 4573
rect 63034 4564 63040 4576
rect 63092 4564 63098 4616
rect 67821 4607 67879 4613
rect 67821 4573 67833 4607
rect 67867 4573 67879 4607
rect 67821 4567 67879 4573
rect 68088 4607 68146 4613
rect 68088 4573 68100 4607
rect 68134 4604 68146 4607
rect 68554 4604 68560 4616
rect 68134 4576 68560 4604
rect 68134 4573 68146 4576
rect 68088 4567 68146 4573
rect 67836 4536 67864 4567
rect 68554 4564 68560 4576
rect 68612 4564 68618 4616
rect 72697 4607 72755 4613
rect 72697 4573 72709 4607
rect 72743 4573 72755 4607
rect 72697 4567 72755 4573
rect 72964 4607 73022 4613
rect 72964 4573 72976 4607
rect 73010 4604 73022 4607
rect 73430 4604 73436 4616
rect 73010 4576 73436 4604
rect 73010 4573 73022 4576
rect 72964 4567 73022 4573
rect 69382 4536 69388 4548
rect 27838 4508 29592 4536
rect 61672 4508 69388 4536
rect 27838 4505 27850 4508
rect 27792 4499 27850 4505
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10965 4471 11023 4477
rect 10965 4468 10977 4471
rect 10284 4440 10977 4468
rect 10284 4428 10290 4440
rect 10965 4437 10977 4440
rect 11011 4437 11023 4471
rect 10965 4431 11023 4437
rect 28166 4428 28172 4480
rect 28224 4468 28230 4480
rect 28626 4468 28632 4480
rect 28224 4440 28632 4468
rect 28224 4428 28230 4440
rect 28626 4428 28632 4440
rect 28684 4468 28690 4480
rect 29564 4477 29592 4508
rect 69382 4496 69388 4508
rect 69440 4536 69446 4548
rect 72712 4536 72740 4567
rect 73430 4564 73436 4576
rect 73488 4564 73494 4616
rect 76929 4607 76987 4613
rect 76929 4573 76941 4607
rect 76975 4573 76987 4607
rect 89456 4604 89484 4635
rect 93946 4604 93952 4616
rect 89456 4576 93808 4604
rect 93907 4576 93952 4604
rect 76929 4567 76987 4573
rect 75914 4536 75920 4548
rect 69440 4508 75920 4536
rect 69440 4496 69446 4508
rect 75914 4496 75920 4508
rect 75972 4496 75978 4548
rect 76469 4539 76527 4545
rect 76469 4505 76481 4539
rect 76515 4536 76527 4539
rect 76742 4536 76748 4548
rect 76515 4508 76748 4536
rect 76515 4505 76527 4508
rect 76469 4499 76527 4505
rect 76742 4496 76748 4508
rect 76800 4496 76806 4548
rect 28905 4471 28963 4477
rect 28905 4468 28917 4471
rect 28684 4440 28917 4468
rect 28684 4428 28690 4440
rect 28905 4437 28917 4440
rect 28951 4437 28963 4471
rect 28905 4431 28963 4437
rect 29549 4471 29607 4477
rect 29549 4437 29561 4471
rect 29595 4437 29607 4471
rect 29549 4431 29607 4437
rect 50154 4428 50160 4480
rect 50212 4468 50218 4480
rect 50525 4471 50583 4477
rect 50525 4468 50537 4471
rect 50212 4440 50537 4468
rect 50212 4428 50218 4440
rect 50525 4437 50537 4440
rect 50571 4437 50583 4471
rect 50525 4431 50583 4437
rect 73890 4428 73896 4480
rect 73948 4468 73954 4480
rect 74077 4471 74135 4477
rect 74077 4468 74089 4471
rect 73948 4440 74089 4468
rect 73948 4428 73954 4440
rect 74077 4437 74089 4440
rect 74123 4468 74135 4471
rect 74442 4468 74448 4480
rect 74123 4440 74448 4468
rect 74123 4437 74135 4440
rect 74077 4431 74135 4437
rect 74442 4428 74448 4440
rect 74500 4468 74506 4480
rect 76944 4468 76972 4567
rect 89708 4539 89766 4545
rect 89708 4505 89720 4539
rect 89754 4536 89766 4539
rect 90358 4536 90364 4548
rect 89754 4508 90364 4536
rect 89754 4505 89766 4508
rect 89708 4499 89766 4505
rect 90358 4496 90364 4508
rect 90416 4496 90422 4548
rect 93780 4536 93808 4576
rect 93946 4564 93952 4576
rect 94004 4564 94010 4616
rect 94133 4607 94191 4613
rect 94133 4573 94145 4607
rect 94179 4604 94191 4607
rect 94682 4604 94688 4616
rect 94179 4576 94688 4604
rect 94179 4573 94191 4576
rect 94133 4567 94191 4573
rect 94682 4564 94688 4576
rect 94740 4564 94746 4616
rect 97353 4607 97411 4613
rect 97353 4573 97365 4607
rect 97399 4604 97411 4607
rect 97460 4604 97488 4712
rect 100294 4700 100300 4712
rect 100352 4700 100358 4752
rect 100772 4740 100800 4768
rect 104897 4743 104955 4749
rect 104897 4740 104909 4743
rect 100772 4712 104909 4740
rect 104897 4709 104909 4712
rect 104943 4740 104955 4743
rect 105078 4740 105084 4752
rect 104943 4712 105084 4740
rect 104943 4709 104955 4712
rect 104897 4703 104955 4709
rect 105078 4700 105084 4712
rect 105136 4700 105142 4752
rect 109954 4700 109960 4752
rect 110012 4740 110018 4752
rect 110012 4712 112576 4740
rect 110012 4700 110018 4712
rect 97626 4672 97632 4684
rect 97587 4644 97632 4672
rect 97626 4632 97632 4644
rect 97684 4632 97690 4684
rect 104989 4675 105047 4681
rect 104989 4641 105001 4675
rect 105035 4672 105047 4675
rect 107838 4672 107844 4684
rect 105035 4644 107844 4672
rect 105035 4641 105047 4644
rect 104989 4635 105047 4641
rect 107838 4632 107844 4644
rect 107896 4632 107902 4684
rect 112438 4672 112444 4684
rect 112399 4644 112444 4672
rect 112438 4632 112444 4644
rect 112496 4632 112502 4684
rect 112548 4681 112576 4712
rect 112533 4675 112591 4681
rect 112533 4641 112545 4675
rect 112579 4641 112591 4675
rect 112533 4635 112591 4641
rect 97399 4576 97488 4604
rect 97537 4607 97595 4613
rect 97399 4573 97411 4576
rect 97353 4567 97411 4573
rect 97537 4573 97549 4607
rect 97583 4573 97595 4607
rect 100202 4604 100208 4616
rect 100163 4576 100208 4604
rect 97537 4567 97595 4573
rect 94038 4536 94044 4548
rect 93780 4508 94044 4536
rect 94038 4496 94044 4508
rect 94096 4496 94102 4548
rect 94314 4536 94320 4548
rect 94275 4508 94320 4536
rect 94314 4496 94320 4508
rect 94372 4496 94378 4548
rect 94590 4496 94596 4548
rect 94648 4536 94654 4548
rect 97552 4536 97580 4567
rect 100202 4564 100208 4576
rect 100260 4564 100266 4616
rect 100389 4607 100447 4613
rect 100389 4573 100401 4607
rect 100435 4604 100447 4607
rect 100938 4604 100944 4616
rect 100435 4576 100944 4604
rect 100435 4573 100447 4576
rect 100389 4567 100447 4573
rect 100938 4564 100944 4576
rect 100996 4564 101002 4616
rect 104710 4604 104716 4616
rect 104671 4576 104716 4604
rect 104710 4564 104716 4576
rect 104768 4564 104774 4616
rect 107378 4604 107384 4616
rect 107339 4576 107384 4604
rect 107378 4564 107384 4576
rect 107436 4564 107442 4616
rect 111337 4607 111395 4613
rect 111337 4573 111349 4607
rect 111383 4604 111395 4607
rect 111383 4576 112024 4604
rect 111383 4573 111395 4576
rect 111337 4567 111395 4573
rect 94648 4508 97580 4536
rect 100220 4536 100248 4564
rect 100478 4536 100484 4548
rect 100220 4508 100484 4536
rect 94648 4496 94654 4508
rect 100478 4496 100484 4508
rect 100536 4496 100542 4548
rect 74500 4440 76972 4468
rect 77113 4471 77171 4477
rect 74500 4428 74506 4440
rect 77113 4437 77125 4471
rect 77159 4468 77171 4471
rect 78582 4468 78588 4480
rect 77159 4440 78588 4468
rect 77159 4437 77171 4440
rect 77113 4431 77171 4437
rect 78582 4428 78588 4440
rect 78640 4428 78646 4480
rect 96798 4428 96804 4480
rect 96856 4468 96862 4480
rect 99006 4468 99012 4480
rect 96856 4440 99012 4468
rect 96856 4428 96862 4440
rect 99006 4428 99012 4440
rect 99064 4468 99070 4480
rect 102318 4468 102324 4480
rect 99064 4440 102324 4468
rect 99064 4428 99070 4440
rect 102318 4428 102324 4440
rect 102376 4468 102382 4480
rect 106458 4468 106464 4480
rect 102376 4440 106464 4468
rect 102376 4428 102382 4440
rect 106458 4428 106464 4440
rect 106516 4468 106522 4480
rect 107010 4468 107016 4480
rect 106516 4440 107016 4468
rect 106516 4428 106522 4440
rect 107010 4428 107016 4440
rect 107068 4428 107074 4480
rect 107194 4468 107200 4480
rect 107155 4440 107200 4468
rect 107194 4428 107200 4440
rect 107252 4428 107258 4480
rect 111150 4468 111156 4480
rect 111111 4440 111156 4468
rect 111150 4428 111156 4440
rect 111208 4428 111214 4480
rect 111996 4477 112024 4576
rect 111981 4471 112039 4477
rect 111981 4437 111993 4471
rect 112027 4437 112039 4471
rect 112346 4468 112352 4480
rect 112307 4440 112352 4468
rect 111981 4431 112039 4437
rect 112346 4428 112352 4440
rect 112404 4428 112410 4480
rect 1104 4378 118864 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 81014 4378
rect 81066 4326 81078 4378
rect 81130 4326 81142 4378
rect 81194 4326 81206 4378
rect 81258 4326 81270 4378
rect 81322 4326 111734 4378
rect 111786 4326 111798 4378
rect 111850 4326 111862 4378
rect 111914 4326 111926 4378
rect 111978 4326 111990 4378
rect 112042 4326 118864 4378
rect 1104 4304 118864 4326
rect 38746 4224 38752 4276
rect 38804 4264 38810 4276
rect 39574 4264 39580 4276
rect 38804 4236 39580 4264
rect 38804 4224 38810 4236
rect 39574 4224 39580 4236
rect 39632 4264 39638 4276
rect 39945 4267 40003 4273
rect 39945 4264 39957 4267
rect 39632 4236 39957 4264
rect 39632 4224 39638 4236
rect 39945 4233 39957 4236
rect 39991 4233 40003 4267
rect 39945 4227 40003 4233
rect 53558 4224 53564 4276
rect 53616 4264 53622 4276
rect 77294 4264 77300 4276
rect 53616 4236 77300 4264
rect 53616 4224 53622 4236
rect 77294 4224 77300 4236
rect 77352 4224 77358 4276
rect 86310 4224 86316 4276
rect 86368 4264 86374 4276
rect 86865 4267 86923 4273
rect 86865 4264 86877 4267
rect 86368 4236 86877 4264
rect 86368 4224 86374 4236
rect 86865 4233 86877 4236
rect 86911 4233 86923 4267
rect 90358 4264 90364 4276
rect 90319 4236 90364 4264
rect 86865 4227 86923 4233
rect 90358 4224 90364 4236
rect 90416 4224 90422 4276
rect 100389 4267 100447 4273
rect 100389 4264 100401 4267
rect 100312 4236 100401 4264
rect 72421 4199 72479 4205
rect 38580 4168 38976 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 2590 4128 2596 4140
rect 1452 4100 2596 4128
rect 1452 4088 1458 4100
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 10226 4128 10232 4140
rect 10187 4100 10232 4128
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4128 10379 4131
rect 10367 4100 16574 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 16546 3992 16574 4100
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 18472 4100 19717 4128
rect 18472 4088 18478 4100
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 19935 4100 22937 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 22925 4097 22937 4100
rect 22971 4128 22983 4131
rect 28353 4131 28411 4137
rect 28353 4128 28365 4131
rect 22971 4100 28365 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 28353 4097 28365 4100
rect 28399 4128 28411 4131
rect 38580 4128 38608 4168
rect 28399 4100 38608 4128
rect 28399 4097 28411 4100
rect 28353 4091 28411 4097
rect 38654 4088 38660 4140
rect 38712 4128 38718 4140
rect 38821 4131 38879 4137
rect 38821 4128 38833 4131
rect 38712 4100 38833 4128
rect 38712 4088 38718 4100
rect 38821 4097 38833 4100
rect 38867 4097 38879 4131
rect 38948 4128 38976 4168
rect 72421 4165 72433 4199
rect 72467 4196 72479 4199
rect 94314 4196 94320 4208
rect 72467 4168 94320 4196
rect 72467 4165 72479 4168
rect 72421 4159 72479 4165
rect 63221 4131 63279 4137
rect 63221 4128 63233 4131
rect 38948 4100 63233 4128
rect 38821 4091 38879 4097
rect 63221 4097 63233 4100
rect 63267 4128 63279 4131
rect 68373 4131 68431 4137
rect 68373 4128 68385 4131
rect 63267 4100 68385 4128
rect 63267 4097 63279 4100
rect 63221 4091 63279 4097
rect 68373 4097 68385 4100
rect 68419 4128 68431 4131
rect 72789 4131 72847 4137
rect 72789 4128 72801 4131
rect 68419 4100 72801 4128
rect 68419 4097 68431 4100
rect 68373 4091 68431 4097
rect 72789 4097 72801 4100
rect 72835 4097 72847 4131
rect 73890 4128 73896 4140
rect 73851 4100 73896 4128
rect 72789 4091 72847 4097
rect 73890 4088 73896 4100
rect 73948 4088 73954 4140
rect 73982 4088 73988 4140
rect 74040 4128 74046 4140
rect 77294 4128 77300 4140
rect 74040 4100 74085 4128
rect 77255 4100 77300 4128
rect 74040 4088 74046 4100
rect 77294 4088 77300 4100
rect 77352 4088 77358 4140
rect 86221 4131 86279 4137
rect 86221 4097 86233 4131
rect 86267 4128 86279 4131
rect 86310 4128 86316 4140
rect 86267 4100 86316 4128
rect 86267 4097 86279 4100
rect 86221 4091 86279 4097
rect 86310 4088 86316 4100
rect 86368 4088 86374 4140
rect 87233 4131 87291 4137
rect 87233 4097 87245 4131
rect 87279 4128 87291 4131
rect 87598 4128 87604 4140
rect 87279 4100 87604 4128
rect 87279 4097 87291 4100
rect 87233 4091 87291 4097
rect 87598 4088 87604 4100
rect 87656 4088 87662 4140
rect 90545 4131 90603 4137
rect 90545 4097 90557 4131
rect 90591 4128 90603 4131
rect 91094 4128 91100 4140
rect 90591 4100 91100 4128
rect 90591 4097 90603 4100
rect 90545 4091 90603 4097
rect 91094 4088 91100 4100
rect 91152 4088 91158 4140
rect 94056 4137 94084 4168
rect 94314 4156 94320 4168
rect 94372 4156 94378 4208
rect 96706 4156 96712 4208
rect 96764 4196 96770 4208
rect 97166 4196 97172 4208
rect 96764 4168 97172 4196
rect 96764 4156 96770 4168
rect 97166 4156 97172 4168
rect 97224 4196 97230 4208
rect 97537 4199 97595 4205
rect 97537 4196 97549 4199
rect 97224 4168 97549 4196
rect 97224 4156 97230 4168
rect 97537 4165 97549 4168
rect 97583 4165 97595 4199
rect 100312 4196 100340 4236
rect 100389 4233 100401 4236
rect 100435 4264 100447 4267
rect 100938 4264 100944 4276
rect 100435 4236 100944 4264
rect 100435 4233 100447 4236
rect 100389 4227 100447 4233
rect 100938 4224 100944 4236
rect 100996 4264 101002 4276
rect 101122 4264 101128 4276
rect 100996 4236 101128 4264
rect 100996 4224 101002 4236
rect 101122 4224 101128 4236
rect 101180 4224 101186 4276
rect 104345 4267 104403 4273
rect 104345 4233 104357 4267
rect 104391 4264 104403 4267
rect 104710 4264 104716 4276
rect 104391 4236 104716 4264
rect 104391 4233 104403 4236
rect 104345 4227 104403 4233
rect 104710 4224 104716 4236
rect 104768 4224 104774 4276
rect 112073 4267 112131 4273
rect 112073 4233 112085 4267
rect 112119 4264 112131 4267
rect 112346 4264 112352 4276
rect 112119 4236 112352 4264
rect 112119 4233 112131 4236
rect 112073 4227 112131 4233
rect 112346 4224 112352 4236
rect 112404 4224 112410 4276
rect 101306 4196 101312 4208
rect 97537 4159 97595 4165
rect 99346 4168 100340 4196
rect 100404 4168 101076 4196
rect 101219 4168 101312 4196
rect 91189 4131 91247 4137
rect 91189 4097 91201 4131
rect 91235 4097 91247 4131
rect 91189 4091 91247 4097
rect 94041 4131 94099 4137
rect 94041 4097 94053 4131
rect 94087 4097 94099 4131
rect 97258 4128 97264 4140
rect 97219 4100 97264 4128
rect 94041 4091 94099 4097
rect 22738 4060 22744 4072
rect 22699 4032 22744 4060
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 28166 4060 28172 4072
rect 28127 4032 28172 4060
rect 28166 4020 28172 4032
rect 28224 4020 28230 4072
rect 38562 4060 38568 4072
rect 38523 4032 38568 4060
rect 38562 4020 38568 4032
rect 38620 4020 38626 4072
rect 45462 4020 45468 4072
rect 45520 4060 45526 4072
rect 50614 4060 50620 4072
rect 45520 4032 50620 4060
rect 45520 4020 45526 4032
rect 50614 4020 50620 4032
rect 50672 4060 50678 4072
rect 59446 4060 59452 4072
rect 50672 4032 59452 4060
rect 50672 4020 50678 4032
rect 59446 4020 59452 4032
rect 59504 4020 59510 4072
rect 63037 4063 63095 4069
rect 63037 4029 63049 4063
rect 63083 4060 63095 4063
rect 63126 4060 63132 4072
rect 63083 4032 63132 4060
rect 63083 4029 63095 4032
rect 63037 4023 63095 4029
rect 63126 4020 63132 4032
rect 63184 4020 63190 4072
rect 68189 4063 68247 4069
rect 68189 4029 68201 4063
rect 68235 4060 68247 4063
rect 69198 4060 69204 4072
rect 68235 4032 69204 4060
rect 68235 4029 68247 4032
rect 68189 4023 68247 4029
rect 69198 4020 69204 4032
rect 69256 4020 69262 4072
rect 74718 4020 74724 4072
rect 74776 4060 74782 4072
rect 77573 4063 77631 4069
rect 77573 4060 77585 4063
rect 74776 4032 77585 4060
rect 74776 4020 74782 4032
rect 77573 4029 77585 4032
rect 77619 4029 77631 4063
rect 86494 4060 86500 4072
rect 86455 4032 86500 4060
rect 77573 4023 77631 4029
rect 35342 3992 35348 4004
rect 16546 3964 35348 3992
rect 35342 3952 35348 3964
rect 35400 3952 35406 4004
rect 68370 3992 68376 4004
rect 39500 3964 68376 3992
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10192 3896 10517 3924
rect 10192 3884 10198 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 20036 3896 20085 3924
rect 20036 3884 20042 3896
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 23109 3927 23167 3933
rect 23109 3893 23121 3927
rect 23155 3924 23167 3927
rect 23750 3924 23756 3936
rect 23155 3896 23756 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 28534 3924 28540 3936
rect 28495 3896 28540 3924
rect 28534 3884 28540 3896
rect 28592 3884 28598 3936
rect 31662 3884 31668 3936
rect 31720 3924 31726 3936
rect 39500 3924 39528 3964
rect 68370 3952 68376 3964
rect 68428 3952 68434 4004
rect 77588 3992 77616 4023
rect 86494 4020 86500 4032
rect 86552 4020 86558 4072
rect 87325 4063 87383 4069
rect 86604 4032 86954 4060
rect 86604 3992 86632 4032
rect 77588 3964 86632 3992
rect 86926 3992 86954 4032
rect 87325 4029 87337 4063
rect 87371 4029 87383 4063
rect 87325 4023 87383 4029
rect 87509 4063 87567 4069
rect 87509 4029 87521 4063
rect 87555 4029 87567 4063
rect 87509 4023 87567 4029
rect 87230 3992 87236 4004
rect 86926 3964 87236 3992
rect 87230 3952 87236 3964
rect 87288 3952 87294 4004
rect 31720 3896 39528 3924
rect 31720 3884 31726 3896
rect 42886 3884 42892 3936
rect 42944 3924 42950 3936
rect 47670 3924 47676 3936
rect 42944 3896 47676 3924
rect 42944 3884 42950 3896
rect 47670 3884 47676 3896
rect 47728 3884 47734 3936
rect 52454 3884 52460 3936
rect 52512 3924 52518 3936
rect 57974 3924 57980 3936
rect 52512 3896 57980 3924
rect 52512 3884 52518 3896
rect 57974 3884 57980 3896
rect 58032 3884 58038 3936
rect 62206 3884 62212 3936
rect 62264 3924 62270 3936
rect 63405 3927 63463 3933
rect 63405 3924 63417 3927
rect 62264 3896 63417 3924
rect 62264 3884 62270 3896
rect 63405 3893 63417 3896
rect 63451 3893 63463 3927
rect 63405 3887 63463 3893
rect 68186 3884 68192 3936
rect 68244 3924 68250 3936
rect 68557 3927 68615 3933
rect 68557 3924 68569 3927
rect 68244 3896 68569 3924
rect 68244 3884 68250 3896
rect 68557 3893 68569 3896
rect 68603 3893 68615 3927
rect 68557 3887 68615 3893
rect 73614 3884 73620 3936
rect 73672 3924 73678 3936
rect 74169 3927 74227 3933
rect 74169 3924 74181 3927
rect 73672 3896 74181 3924
rect 73672 3884 73678 3896
rect 74169 3893 74181 3896
rect 74215 3893 74227 3927
rect 74169 3887 74227 3893
rect 86037 3927 86095 3933
rect 86037 3893 86049 3927
rect 86083 3924 86095 3927
rect 86310 3924 86316 3936
rect 86083 3896 86316 3924
rect 86083 3893 86095 3896
rect 86037 3887 86095 3893
rect 86310 3884 86316 3896
rect 86368 3884 86374 3936
rect 86494 3884 86500 3936
rect 86552 3924 86558 3936
rect 87340 3924 87368 4023
rect 87524 3992 87552 4023
rect 90726 4020 90732 4072
rect 90784 4060 90790 4072
rect 91204 4060 91232 4091
rect 97258 4088 97264 4100
rect 97316 4088 97322 4140
rect 99346 4128 99374 4168
rect 97368 4100 99374 4128
rect 100205 4131 100263 4137
rect 90784 4032 91232 4060
rect 90784 4020 90790 4032
rect 93854 4020 93860 4072
rect 93912 4060 93918 4072
rect 94317 4063 94375 4069
rect 94317 4060 94329 4063
rect 93912 4032 94329 4060
rect 93912 4020 93918 4032
rect 94317 4029 94329 4032
rect 94363 4060 94375 4063
rect 94590 4060 94596 4072
rect 94363 4032 94596 4060
rect 94363 4029 94375 4032
rect 94317 4023 94375 4029
rect 94590 4020 94596 4032
rect 94648 4020 94654 4072
rect 94682 4020 94688 4072
rect 94740 4060 94746 4072
rect 97368 4060 97396 4100
rect 100205 4097 100217 4131
rect 100251 4128 100263 4131
rect 100404 4128 100432 4168
rect 100251 4100 100432 4128
rect 100251 4097 100263 4100
rect 100205 4091 100263 4097
rect 100478 4088 100484 4140
rect 100536 4128 100542 4140
rect 100941 4131 100999 4137
rect 100941 4128 100953 4131
rect 100536 4100 100953 4128
rect 100536 4088 100542 4100
rect 100941 4097 100953 4100
rect 100987 4097 100999 4131
rect 100941 4091 100999 4097
rect 94740 4032 97396 4060
rect 100021 4063 100079 4069
rect 94740 4020 94746 4032
rect 100021 4029 100033 4063
rect 100067 4060 100079 4063
rect 100386 4060 100392 4072
rect 100067 4032 100392 4060
rect 100067 4029 100079 4032
rect 100021 4023 100079 4029
rect 100386 4020 100392 4032
rect 100444 4060 100450 4072
rect 101048 4060 101076 4168
rect 101306 4156 101312 4168
rect 101364 4196 101370 4208
rect 101364 4168 101904 4196
rect 101364 4156 101370 4168
rect 101122 4088 101128 4140
rect 101180 4128 101186 4140
rect 101490 4128 101496 4140
rect 101180 4100 101225 4128
rect 101451 4100 101496 4128
rect 101180 4088 101186 4100
rect 101490 4088 101496 4100
rect 101548 4088 101554 4140
rect 101766 4128 101772 4140
rect 101727 4100 101772 4128
rect 101766 4088 101772 4100
rect 101824 4088 101830 4140
rect 101876 4128 101904 4168
rect 104820 4168 105216 4196
rect 104253 4131 104311 4137
rect 104253 4128 104265 4131
rect 101876 4100 104265 4128
rect 104253 4097 104265 4100
rect 104299 4097 104311 4131
rect 104253 4091 104311 4097
rect 104437 4131 104495 4137
rect 104437 4097 104449 4131
rect 104483 4128 104495 4131
rect 104820 4128 104848 4168
rect 104483 4100 104848 4128
rect 104897 4131 104955 4137
rect 104483 4097 104495 4100
rect 104437 4091 104495 4097
rect 104897 4097 104909 4131
rect 104943 4097 104955 4131
rect 105078 4128 105084 4140
rect 105039 4100 105084 4128
rect 104897 4091 104955 4097
rect 101674 4060 101680 4072
rect 100444 4032 100984 4060
rect 101048 4032 101680 4060
rect 100444 4020 100450 4032
rect 87524 3964 91600 3992
rect 86552 3896 87368 3924
rect 86552 3884 86558 3896
rect 89070 3884 89076 3936
rect 89128 3924 89134 3936
rect 89349 3927 89407 3933
rect 89349 3924 89361 3927
rect 89128 3896 89361 3924
rect 89128 3884 89134 3896
rect 89349 3893 89361 3896
rect 89395 3893 89407 3927
rect 89349 3887 89407 3893
rect 90542 3884 90548 3936
rect 90600 3924 90606 3936
rect 91005 3927 91063 3933
rect 91005 3924 91017 3927
rect 90600 3896 91017 3924
rect 90600 3884 90606 3896
rect 91005 3893 91017 3896
rect 91051 3893 91063 3927
rect 91572 3924 91600 3964
rect 91646 3952 91652 4004
rect 91704 3992 91710 4004
rect 100956 3992 100984 4032
rect 101674 4020 101680 4032
rect 101732 4060 101738 4072
rect 104452 4060 104480 4091
rect 101732 4032 104480 4060
rect 101732 4020 101738 4032
rect 104912 3992 104940 4091
rect 105078 4088 105084 4100
rect 105136 4088 105142 4140
rect 105188 4128 105216 4168
rect 107194 4156 107200 4208
rect 107252 4196 107258 4208
rect 107350 4199 107408 4205
rect 107350 4196 107362 4199
rect 107252 4168 107362 4196
rect 107252 4156 107258 4168
rect 107350 4165 107362 4168
rect 107396 4165 107408 4199
rect 107350 4159 107408 4165
rect 110960 4199 111018 4205
rect 110960 4165 110972 4199
rect 111006 4196 111018 4199
rect 111150 4196 111156 4208
rect 111006 4168 111156 4196
rect 111006 4165 111018 4168
rect 110960 4159 111018 4165
rect 111150 4156 111156 4168
rect 111208 4156 111214 4208
rect 117958 4196 117964 4208
rect 117919 4168 117964 4196
rect 117958 4156 117964 4168
rect 118016 4156 118022 4208
rect 118145 4131 118203 4137
rect 118145 4128 118157 4131
rect 105188 4100 108160 4128
rect 107102 4060 107108 4072
rect 107063 4032 107108 4060
rect 107102 4020 107108 4032
rect 107160 4020 107166 4072
rect 108132 4060 108160 4100
rect 109144 4100 118157 4128
rect 109144 4060 109172 4100
rect 118145 4097 118157 4100
rect 118191 4097 118203 4131
rect 118145 4091 118203 4097
rect 108132 4032 109172 4060
rect 110693 4063 110751 4069
rect 110693 4029 110705 4063
rect 110739 4029 110751 4063
rect 110693 4023 110751 4029
rect 109678 3992 109684 4004
rect 91704 3964 99374 3992
rect 100956 3964 104940 3992
rect 108040 3964 109684 3992
rect 91704 3952 91710 3964
rect 97994 3924 98000 3936
rect 91572 3896 98000 3924
rect 91005 3887 91063 3893
rect 97994 3884 98000 3896
rect 98052 3884 98058 3936
rect 99346 3924 99374 3964
rect 103606 3924 103612 3936
rect 99346 3896 103612 3924
rect 103606 3884 103612 3896
rect 103664 3884 103670 3936
rect 104894 3924 104900 3936
rect 104855 3896 104900 3924
rect 104894 3884 104900 3896
rect 104952 3884 104958 3936
rect 105170 3884 105176 3936
rect 105228 3924 105234 3936
rect 108040 3924 108068 3964
rect 109678 3952 109684 3964
rect 109736 3952 109742 4004
rect 108482 3924 108488 3936
rect 105228 3896 108068 3924
rect 108443 3896 108488 3924
rect 105228 3884 105234 3896
rect 108482 3884 108488 3896
rect 108540 3884 108546 3936
rect 110708 3924 110736 4023
rect 110966 3924 110972 3936
rect 110708 3896 110972 3924
rect 110966 3884 110972 3896
rect 111024 3884 111030 3936
rect 1104 3834 118864 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 118864 3834
rect 1104 3760 118864 3782
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 59262 3720 59268 3732
rect 2924 3692 55904 3720
rect 59223 3692 59268 3720
rect 2924 3680 2930 3692
rect 35342 3612 35348 3664
rect 35400 3652 35406 3664
rect 38378 3652 38384 3664
rect 35400 3624 38384 3652
rect 35400 3612 35406 3624
rect 38378 3612 38384 3624
rect 38436 3652 38442 3664
rect 45462 3652 45468 3664
rect 38436 3624 45468 3652
rect 38436 3612 38442 3624
rect 45462 3612 45468 3624
rect 45520 3612 45526 3664
rect 45646 3652 45652 3664
rect 45607 3624 45652 3652
rect 45646 3612 45652 3624
rect 45704 3612 45710 3664
rect 46477 3655 46535 3661
rect 46477 3621 46489 3655
rect 46523 3652 46535 3655
rect 47578 3652 47584 3664
rect 46523 3624 47584 3652
rect 46523 3621 46535 3624
rect 46477 3615 46535 3621
rect 47578 3612 47584 3624
rect 47636 3612 47642 3664
rect 47670 3612 47676 3664
rect 47728 3652 47734 3664
rect 52454 3652 52460 3664
rect 47728 3624 52460 3652
rect 47728 3612 47734 3624
rect 52454 3612 52460 3624
rect 52512 3612 52518 3664
rect 55876 3652 55904 3692
rect 59262 3680 59268 3692
rect 59320 3680 59326 3732
rect 79134 3720 79140 3732
rect 59372 3692 79140 3720
rect 59372 3652 59400 3692
rect 79134 3680 79140 3692
rect 79192 3680 79198 3732
rect 83737 3723 83795 3729
rect 83737 3689 83749 3723
rect 83783 3720 83795 3723
rect 83783 3692 87184 3720
rect 83783 3689 83795 3692
rect 83737 3683 83795 3689
rect 52564 3624 54248 3652
rect 55876 3624 59400 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 52564 3584 52592 3624
rect 52730 3584 52736 3596
rect 1728 3556 52592 3584
rect 52691 3556 52736 3584
rect 1728 3544 1734 3556
rect 52730 3544 52736 3556
rect 52788 3544 52794 3596
rect 54110 3584 54116 3596
rect 54071 3556 54116 3584
rect 54110 3544 54116 3556
rect 54168 3544 54174 3596
rect 54220 3584 54248 3624
rect 59446 3612 59452 3664
rect 59504 3652 59510 3664
rect 73982 3652 73988 3664
rect 59504 3624 73988 3652
rect 59504 3612 59510 3624
rect 73982 3612 73988 3624
rect 74040 3612 74046 3664
rect 87156 3652 87184 3692
rect 87230 3680 87236 3732
rect 87288 3720 87294 3732
rect 91554 3720 91560 3732
rect 87288 3692 91560 3720
rect 87288 3680 87294 3692
rect 91554 3680 91560 3692
rect 91612 3680 91618 3732
rect 91738 3720 91744 3732
rect 91699 3692 91744 3720
rect 91738 3680 91744 3692
rect 91796 3680 91802 3732
rect 92474 3720 92480 3732
rect 92435 3692 92480 3720
rect 92474 3680 92480 3692
rect 92532 3680 92538 3732
rect 97994 3720 98000 3732
rect 97955 3692 98000 3720
rect 97994 3680 98000 3692
rect 98052 3680 98058 3732
rect 100113 3723 100171 3729
rect 100113 3689 100125 3723
rect 100159 3720 100171 3723
rect 100294 3720 100300 3732
rect 100159 3692 100300 3720
rect 100159 3689 100171 3692
rect 100113 3683 100171 3689
rect 100294 3680 100300 3692
rect 100352 3680 100358 3732
rect 107289 3723 107347 3729
rect 107289 3689 107301 3723
rect 107335 3720 107347 3723
rect 107378 3720 107384 3732
rect 107335 3692 107384 3720
rect 107335 3689 107347 3692
rect 107289 3683 107347 3689
rect 107378 3680 107384 3692
rect 107436 3680 107442 3732
rect 109770 3680 109776 3732
rect 109828 3720 109834 3732
rect 112257 3723 112315 3729
rect 112257 3720 112269 3723
rect 109828 3692 112269 3720
rect 109828 3680 109834 3692
rect 112257 3689 112269 3692
rect 112303 3689 112315 3723
rect 117498 3720 117504 3732
rect 112257 3683 112315 3689
rect 113146 3692 117504 3720
rect 92201 3655 92259 3661
rect 92201 3652 92213 3655
rect 87156 3624 92213 3652
rect 92201 3621 92213 3624
rect 92247 3621 92259 3655
rect 92201 3615 92259 3621
rect 94317 3655 94375 3661
rect 94317 3621 94329 3655
rect 94363 3652 94375 3655
rect 94682 3652 94688 3664
rect 94363 3624 94688 3652
rect 94363 3621 94375 3624
rect 94317 3615 94375 3621
rect 94682 3612 94688 3624
rect 94740 3612 94746 3664
rect 99101 3655 99159 3661
rect 99101 3621 99113 3655
rect 99147 3652 99159 3655
rect 113146 3652 113174 3692
rect 117498 3680 117504 3692
rect 117556 3680 117562 3732
rect 99147 3624 113174 3652
rect 99147 3621 99159 3624
rect 99101 3615 99159 3621
rect 56137 3587 56195 3593
rect 56137 3584 56149 3587
rect 54220 3556 56149 3584
rect 56137 3553 56149 3556
rect 56183 3553 56195 3587
rect 64322 3584 64328 3596
rect 56137 3547 56195 3553
rect 57072 3556 60734 3584
rect 64283 3556 64328 3584
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 2406 3516 2412 3528
rect 2367 3488 2412 3516
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 2590 3476 2596 3528
rect 2648 3516 2654 3528
rect 10134 3516 10140 3528
rect 2648 3488 6914 3516
rect 10095 3488 10140 3516
rect 2648 3476 2654 3488
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2869 3451 2927 3457
rect 2869 3448 2881 3451
rect 2004 3420 2881 3448
rect 2004 3408 2010 3420
rect 2869 3417 2881 3420
rect 2915 3417 2927 3451
rect 6886 3448 6914 3488
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 19978 3516 19984 3528
rect 19939 3488 19984 3516
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 23750 3516 23756 3528
rect 23711 3488 23756 3516
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 28534 3516 28540 3528
rect 28495 3488 28540 3516
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 38470 3516 38476 3528
rect 28966 3488 37964 3516
rect 38431 3488 38476 3516
rect 28966 3448 28994 3488
rect 6886 3420 28994 3448
rect 37645 3451 37703 3457
rect 2869 3411 2927 3417
rect 37645 3417 37657 3451
rect 37691 3417 37703 3451
rect 37826 3448 37832 3460
rect 37787 3420 37832 3448
rect 37645 3411 37703 3417
rect 382 3340 388 3392
rect 440 3380 446 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 440 3352 1593 3380
rect 440 3340 446 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 1581 3343 1639 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 9953 3383 10011 3389
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 10042 3380 10048 3392
rect 9999 3352 10048 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19797 3383 19855 3389
rect 19797 3380 19809 3383
rect 19484 3352 19809 3380
rect 19484 3340 19490 3352
rect 19797 3349 19809 3352
rect 19843 3349 19855 3383
rect 19797 3343 19855 3349
rect 23569 3383 23627 3389
rect 23569 3349 23581 3383
rect 23615 3380 23627 3383
rect 24394 3380 24400 3392
rect 23615 3352 24400 3380
rect 23615 3349 23627 3352
rect 23569 3343 23627 3349
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 28353 3383 28411 3389
rect 28353 3349 28365 3383
rect 28399 3380 28411 3383
rect 28442 3380 28448 3392
rect 28399 3352 28448 3380
rect 28399 3349 28411 3352
rect 28353 3343 28411 3349
rect 28442 3340 28448 3352
rect 28500 3340 28506 3392
rect 37660 3380 37688 3411
rect 37826 3408 37832 3420
rect 37884 3408 37890 3460
rect 37936 3448 37964 3488
rect 38470 3476 38476 3488
rect 38528 3476 38534 3528
rect 38562 3476 38568 3528
rect 38620 3525 38626 3528
rect 38620 3519 38643 3525
rect 38631 3485 38643 3519
rect 42886 3516 42892 3528
rect 38620 3479 38643 3485
rect 38672 3488 42892 3516
rect 38620 3476 38626 3479
rect 38672 3448 38700 3488
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 45462 3476 45468 3528
rect 45520 3516 45526 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 45520 3488 45565 3516
rect 46216 3488 46305 3516
rect 45520 3476 45526 3488
rect 37936 3420 38700 3448
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 46106 3448 46112 3460
rect 40736 3420 46112 3448
rect 40736 3408 40742 3420
rect 46106 3408 46112 3420
rect 46164 3408 46170 3460
rect 38749 3383 38807 3389
rect 38749 3380 38761 3383
rect 37660 3352 38761 3380
rect 38749 3349 38761 3352
rect 38795 3349 38807 3383
rect 38749 3343 38807 3349
rect 40218 3340 40224 3392
rect 40276 3380 40282 3392
rect 46216 3380 46244 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 46474 3476 46480 3528
rect 46532 3516 46538 3528
rect 47397 3519 47455 3525
rect 47397 3516 47409 3519
rect 46532 3488 47409 3516
rect 46532 3476 46538 3488
rect 47397 3485 47409 3488
rect 47443 3485 47455 3519
rect 47578 3516 47584 3528
rect 47539 3488 47584 3516
rect 47397 3479 47455 3485
rect 47578 3476 47584 3488
rect 47636 3476 47642 3528
rect 50154 3516 50160 3528
rect 50115 3488 50160 3516
rect 50154 3476 50160 3488
rect 50212 3476 50218 3528
rect 52454 3516 52460 3528
rect 52415 3488 52460 3516
rect 52454 3476 52460 3488
rect 52512 3476 52518 3528
rect 52822 3476 52828 3528
rect 52880 3516 52886 3528
rect 55953 3519 56011 3525
rect 52880 3488 53512 3516
rect 52880 3476 52886 3488
rect 47765 3451 47823 3457
rect 47765 3417 47777 3451
rect 47811 3448 47823 3451
rect 47811 3420 51074 3448
rect 47811 3417 47823 3420
rect 47765 3411 47823 3417
rect 40276 3352 46244 3380
rect 40276 3340 40282 3352
rect 46382 3340 46388 3392
rect 46440 3380 46446 3392
rect 50341 3383 50399 3389
rect 50341 3380 50353 3383
rect 46440 3352 50353 3380
rect 46440 3340 46446 3352
rect 50341 3349 50353 3352
rect 50387 3349 50399 3383
rect 51046 3380 51074 3420
rect 53282 3408 53288 3460
rect 53340 3448 53346 3460
rect 53377 3451 53435 3457
rect 53377 3448 53389 3451
rect 53340 3420 53389 3448
rect 53340 3408 53346 3420
rect 53377 3417 53389 3420
rect 53423 3417 53435 3451
rect 53484 3448 53512 3488
rect 55953 3485 55965 3519
rect 55999 3516 56011 3519
rect 56962 3516 56968 3528
rect 55999 3488 56968 3516
rect 55999 3485 56011 3488
rect 55953 3479 56011 3485
rect 56962 3476 56968 3488
rect 57020 3476 57026 3528
rect 57072 3448 57100 3556
rect 59081 3519 59139 3525
rect 59081 3485 59093 3519
rect 59127 3485 59139 3519
rect 59081 3479 59139 3485
rect 53484 3420 57100 3448
rect 53377 3411 53435 3417
rect 59096 3380 59124 3479
rect 60706 3448 60734 3556
rect 64322 3544 64328 3556
rect 64380 3544 64386 3596
rect 78582 3544 78588 3596
rect 78640 3584 78646 3596
rect 83645 3587 83703 3593
rect 83645 3584 83657 3587
rect 78640 3556 83657 3584
rect 78640 3544 78646 3556
rect 83645 3553 83657 3556
rect 83691 3553 83703 3587
rect 86218 3584 86224 3596
rect 86179 3556 86224 3584
rect 83645 3547 83703 3553
rect 86218 3544 86224 3556
rect 86276 3544 86282 3596
rect 87598 3584 87604 3596
rect 87511 3556 87604 3584
rect 87598 3544 87604 3556
rect 87656 3584 87662 3596
rect 91738 3584 91744 3596
rect 87656 3556 91744 3584
rect 87656 3544 87662 3556
rect 91738 3544 91744 3556
rect 91796 3544 91802 3596
rect 91922 3584 91928 3596
rect 91883 3556 91928 3584
rect 91922 3544 91928 3556
rect 91980 3544 91986 3596
rect 93946 3584 93952 3596
rect 93907 3556 93952 3584
rect 93946 3544 93952 3556
rect 94004 3544 94010 3596
rect 97166 3584 97172 3596
rect 97127 3556 97172 3584
rect 97166 3544 97172 3556
rect 97224 3544 97230 3596
rect 101306 3584 101312 3596
rect 100128 3556 101312 3584
rect 62206 3516 62212 3528
rect 62167 3488 62212 3516
rect 62206 3476 62212 3488
rect 62264 3476 62270 3528
rect 64046 3516 64052 3528
rect 64007 3488 64052 3516
rect 64046 3476 64052 3488
rect 64104 3476 64110 3528
rect 66073 3519 66131 3525
rect 66073 3485 66085 3519
rect 66119 3516 66131 3519
rect 66806 3516 66812 3528
rect 66119 3488 66812 3516
rect 66119 3485 66131 3488
rect 66073 3479 66131 3485
rect 66806 3476 66812 3488
rect 66864 3476 66870 3528
rect 67821 3519 67879 3525
rect 67821 3485 67833 3519
rect 67867 3516 67879 3519
rect 68830 3516 68836 3528
rect 67867 3488 68836 3516
rect 67867 3485 67879 3488
rect 67821 3479 67879 3485
rect 68830 3476 68836 3488
rect 68888 3476 68894 3528
rect 73890 3476 73896 3528
rect 73948 3516 73954 3528
rect 74169 3519 74227 3525
rect 74169 3516 74181 3519
rect 73948 3488 74181 3516
rect 73948 3476 73954 3488
rect 74169 3485 74181 3488
rect 74215 3485 74227 3519
rect 83550 3516 83556 3528
rect 83511 3488 83556 3516
rect 74169 3479 74227 3485
rect 83550 3476 83556 3488
rect 83608 3476 83614 3528
rect 86310 3476 86316 3528
rect 86368 3516 86374 3528
rect 86477 3519 86535 3525
rect 86477 3516 86489 3519
rect 86368 3488 86489 3516
rect 86368 3476 86374 3488
rect 86477 3485 86489 3488
rect 86523 3485 86535 3519
rect 86477 3479 86535 3485
rect 66441 3451 66499 3457
rect 66441 3448 66453 3451
rect 60706 3420 66453 3448
rect 66441 3417 66453 3420
rect 66487 3417 66499 3451
rect 66441 3411 66499 3417
rect 68189 3451 68247 3457
rect 68189 3417 68201 3451
rect 68235 3417 68247 3451
rect 68189 3411 68247 3417
rect 51046 3352 59124 3380
rect 50341 3343 50399 3349
rect 61746 3340 61752 3392
rect 61804 3380 61810 3392
rect 62301 3383 62359 3389
rect 62301 3380 62313 3383
rect 61804 3352 62313 3380
rect 61804 3340 61810 3352
rect 62301 3349 62313 3352
rect 62347 3349 62359 3383
rect 62301 3343 62359 3349
rect 62390 3340 62396 3392
rect 62448 3380 62454 3392
rect 68204 3380 68232 3411
rect 62448 3352 68232 3380
rect 73985 3383 74043 3389
rect 62448 3340 62454 3352
rect 73985 3349 73997 3383
rect 74031 3380 74043 3383
rect 74534 3380 74540 3392
rect 74031 3352 74540 3380
rect 74031 3349 74043 3352
rect 73985 3343 74043 3349
rect 74534 3340 74540 3352
rect 74592 3340 74598 3392
rect 83642 3340 83648 3392
rect 83700 3380 83706 3392
rect 87616 3389 87644 3544
rect 88702 3516 88708 3528
rect 88663 3488 88708 3516
rect 88702 3476 88708 3488
rect 88760 3516 88766 3528
rect 89073 3519 89131 3525
rect 89073 3516 89085 3519
rect 88760 3488 89085 3516
rect 88760 3476 88766 3488
rect 89073 3485 89085 3488
rect 89119 3516 89131 3519
rect 89441 3519 89499 3525
rect 89441 3516 89453 3519
rect 89119 3488 89453 3516
rect 89119 3485 89131 3488
rect 89073 3479 89131 3485
rect 89441 3485 89453 3488
rect 89487 3516 89499 3519
rect 89993 3519 90051 3525
rect 89487 3488 89714 3516
rect 89487 3485 89499 3488
rect 89441 3479 89499 3485
rect 87690 3408 87696 3460
rect 87748 3448 87754 3460
rect 89686 3448 89714 3488
rect 89993 3485 90005 3519
rect 90039 3516 90051 3519
rect 91646 3516 91652 3528
rect 90039 3488 91652 3516
rect 90039 3485 90051 3488
rect 89993 3479 90051 3485
rect 91646 3476 91652 3488
rect 91704 3476 91710 3528
rect 92057 3519 92115 3525
rect 92057 3485 92069 3519
rect 92103 3516 92115 3519
rect 95050 3516 95056 3528
rect 92103 3488 95056 3516
rect 92103 3485 92115 3488
rect 92057 3479 92115 3485
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 95145 3519 95203 3525
rect 95145 3485 95157 3519
rect 95191 3516 95203 3519
rect 97077 3519 97135 3525
rect 95191 3488 96660 3516
rect 95191 3485 95203 3488
rect 95145 3479 95203 3485
rect 90637 3451 90695 3457
rect 90637 3448 90649 3451
rect 87748 3420 89576 3448
rect 89686 3420 90649 3448
rect 87748 3408 87754 3420
rect 83921 3383 83979 3389
rect 83921 3380 83933 3383
rect 83700 3352 83933 3380
rect 83700 3340 83706 3352
rect 83921 3349 83933 3352
rect 83967 3349 83979 3383
rect 83921 3343 83979 3349
rect 87601 3383 87659 3389
rect 87601 3349 87613 3383
rect 87647 3349 87659 3383
rect 89548 3380 89576 3420
rect 90637 3417 90649 3420
rect 90683 3448 90695 3451
rect 91557 3451 91615 3457
rect 91557 3448 91569 3451
rect 90683 3420 91569 3448
rect 90683 3417 90695 3420
rect 90637 3411 90695 3417
rect 91557 3417 91569 3420
rect 91603 3417 91615 3451
rect 91738 3448 91744 3460
rect 91699 3420 91744 3448
rect 91557 3411 91615 3417
rect 91738 3408 91744 3420
rect 91796 3408 91802 3460
rect 91830 3408 91836 3460
rect 91888 3448 91894 3460
rect 92385 3451 92443 3457
rect 92385 3448 92397 3451
rect 91888 3420 92397 3448
rect 91888 3408 91894 3420
rect 92385 3417 92397 3420
rect 92431 3417 92443 3451
rect 92385 3411 92443 3417
rect 89622 3380 89628 3392
rect 89548 3352 89628 3380
rect 87601 3343 87659 3349
rect 89622 3340 89628 3352
rect 89680 3340 89686 3392
rect 91186 3340 91192 3392
rect 91244 3380 91250 3392
rect 94409 3383 94467 3389
rect 94409 3380 94421 3383
rect 91244 3352 94421 3380
rect 91244 3340 91250 3352
rect 94409 3349 94421 3352
rect 94455 3349 94467 3383
rect 94958 3380 94964 3392
rect 94919 3352 94964 3380
rect 94409 3343 94467 3349
rect 94958 3340 94964 3352
rect 95016 3340 95022 3392
rect 96632 3389 96660 3488
rect 97077 3485 97089 3519
rect 97123 3516 97135 3519
rect 99282 3516 99288 3528
rect 97123 3488 99288 3516
rect 97123 3485 97135 3488
rect 97077 3479 97135 3485
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 100128 3525 100156 3556
rect 101306 3544 101312 3556
rect 101364 3544 101370 3596
rect 101674 3584 101680 3596
rect 101635 3556 101680 3584
rect 101674 3544 101680 3556
rect 101732 3544 101738 3596
rect 101766 3544 101772 3596
rect 101824 3584 101830 3596
rect 102162 3587 102220 3593
rect 102162 3584 102174 3587
rect 101824 3556 102174 3584
rect 101824 3544 101830 3556
rect 102162 3553 102174 3556
rect 102208 3553 102220 3587
rect 102162 3547 102220 3553
rect 103606 3544 103612 3596
rect 103664 3584 103670 3596
rect 107841 3587 107899 3593
rect 107841 3584 107853 3587
rect 103664 3556 107853 3584
rect 103664 3544 103670 3556
rect 107841 3553 107853 3556
rect 107887 3553 107899 3587
rect 108482 3584 108488 3596
rect 107841 3547 107899 3553
rect 108316 3556 108488 3584
rect 100113 3519 100171 3525
rect 100113 3485 100125 3519
rect 100159 3485 100171 3519
rect 100113 3479 100171 3485
rect 100297 3519 100355 3525
rect 100297 3485 100309 3519
rect 100343 3516 100355 3519
rect 100386 3516 100392 3528
rect 100343 3488 100392 3516
rect 100343 3485 100355 3488
rect 100297 3479 100355 3485
rect 100386 3476 100392 3488
rect 100444 3476 100450 3528
rect 101490 3476 101496 3528
rect 101548 3516 101554 3528
rect 102045 3519 102103 3525
rect 102045 3516 102057 3519
rect 101548 3488 102057 3516
rect 101548 3476 101554 3488
rect 102045 3485 102057 3488
rect 102091 3516 102103 3519
rect 107657 3519 107715 3525
rect 102091 3488 104204 3516
rect 102091 3485 102103 3488
rect 102045 3479 102103 3485
rect 97258 3408 97264 3460
rect 97316 3448 97322 3460
rect 97905 3451 97963 3457
rect 97905 3448 97917 3451
rect 97316 3420 97917 3448
rect 97316 3408 97322 3420
rect 97905 3417 97917 3420
rect 97951 3448 97963 3451
rect 97951 3420 98132 3448
rect 97951 3417 97963 3420
rect 97905 3411 97963 3417
rect 96617 3383 96675 3389
rect 96617 3349 96629 3383
rect 96663 3349 96675 3383
rect 96982 3380 96988 3392
rect 96943 3352 96988 3380
rect 96617 3343 96675 3349
rect 96982 3340 96988 3352
rect 97040 3340 97046 3392
rect 98104 3380 98132 3420
rect 98178 3408 98184 3460
rect 98236 3448 98242 3460
rect 98825 3451 98883 3457
rect 98825 3448 98837 3451
rect 98236 3420 98837 3448
rect 98236 3408 98242 3420
rect 98825 3417 98837 3420
rect 98871 3417 98883 3451
rect 104176 3448 104204 3488
rect 107657 3485 107669 3519
rect 107703 3516 107715 3519
rect 108316 3516 108344 3556
rect 108482 3544 108488 3556
rect 108540 3584 108546 3596
rect 112349 3587 112407 3593
rect 112349 3584 112361 3587
rect 108540 3556 112361 3584
rect 108540 3544 108546 3556
rect 112349 3553 112361 3556
rect 112395 3553 112407 3587
rect 112349 3547 112407 3553
rect 107703 3488 108344 3516
rect 107703 3485 107715 3488
rect 107657 3479 107715 3485
rect 108390 3476 108396 3528
rect 108448 3516 108454 3528
rect 108669 3519 108727 3525
rect 108669 3516 108681 3519
rect 108448 3488 108681 3516
rect 108448 3476 108454 3488
rect 108669 3485 108681 3488
rect 108715 3485 108727 3519
rect 108669 3479 108727 3485
rect 112128 3519 112186 3525
rect 112128 3485 112140 3519
rect 112174 3516 112186 3519
rect 115566 3516 115572 3528
rect 112174 3485 112208 3516
rect 112128 3479 112208 3485
rect 111978 3448 111984 3460
rect 98825 3411 98883 3417
rect 99346 3420 102364 3448
rect 104176 3420 109034 3448
rect 111939 3420 111984 3448
rect 99346 3380 99374 3420
rect 98104 3352 99374 3380
rect 100754 3340 100760 3392
rect 100812 3380 100818 3392
rect 102336 3389 102364 3420
rect 101953 3383 102011 3389
rect 101953 3380 101965 3383
rect 100812 3352 101965 3380
rect 100812 3340 100818 3352
rect 101953 3349 101965 3352
rect 101999 3349 102011 3383
rect 101953 3343 102011 3349
rect 102321 3383 102379 3389
rect 102321 3349 102333 3383
rect 102367 3349 102379 3383
rect 102321 3343 102379 3349
rect 107749 3383 107807 3389
rect 107749 3349 107761 3383
rect 107795 3380 107807 3383
rect 108485 3383 108543 3389
rect 108485 3380 108497 3383
rect 107795 3352 108497 3380
rect 107795 3349 107807 3352
rect 107749 3343 107807 3349
rect 108485 3349 108497 3352
rect 108531 3349 108543 3383
rect 109006 3380 109034 3420
rect 111978 3408 111984 3420
rect 112036 3408 112042 3460
rect 112180 3448 112208 3479
rect 112456 3488 115572 3516
rect 112346 3448 112352 3460
rect 112180 3420 112352 3448
rect 112346 3408 112352 3420
rect 112404 3408 112410 3460
rect 112456 3380 112484 3488
rect 115566 3476 115572 3488
rect 115624 3476 115630 3528
rect 117406 3476 117412 3528
rect 117464 3516 117470 3528
rect 117869 3519 117927 3525
rect 117869 3516 117881 3519
rect 117464 3488 117881 3516
rect 117464 3476 117470 3488
rect 117869 3485 117881 3488
rect 117915 3485 117927 3519
rect 117869 3479 117927 3485
rect 112622 3380 112628 3392
rect 109006 3352 112484 3380
rect 112583 3352 112628 3380
rect 108485 3343 108543 3349
rect 112622 3340 112628 3352
rect 112680 3340 112686 3392
rect 118053 3383 118111 3389
rect 118053 3349 118065 3383
rect 118099 3380 118111 3383
rect 118142 3380 118148 3392
rect 118099 3352 118148 3380
rect 118099 3349 118111 3352
rect 118053 3343 118111 3349
rect 118142 3340 118148 3352
rect 118200 3340 118206 3392
rect 1104 3290 118864 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 81014 3290
rect 81066 3238 81078 3290
rect 81130 3238 81142 3290
rect 81194 3238 81206 3290
rect 81258 3238 81270 3290
rect 81322 3238 111734 3290
rect 111786 3238 111798 3290
rect 111850 3238 111862 3290
rect 111914 3238 111926 3290
rect 111978 3238 111990 3290
rect 112042 3238 118864 3290
rect 1104 3216 118864 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 1452 3148 2237 3176
rect 1452 3136 1458 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 6886 3148 45968 3176
rect 1486 3068 1492 3120
rect 1544 3108 1550 3120
rect 6886 3108 6914 3148
rect 45940 3108 45968 3148
rect 46198 3136 46204 3188
rect 46256 3176 46262 3188
rect 51902 3176 51908 3188
rect 46256 3148 51908 3176
rect 46256 3136 46262 3148
rect 51902 3136 51908 3148
rect 51960 3136 51966 3188
rect 51997 3179 52055 3185
rect 51997 3145 52009 3179
rect 52043 3176 52055 3179
rect 53282 3176 53288 3188
rect 52043 3148 52960 3176
rect 53243 3148 53288 3176
rect 52043 3145 52055 3148
rect 51997 3139 52055 3145
rect 52822 3108 52828 3120
rect 1544 3080 6914 3108
rect 16546 3080 43484 3108
rect 45940 3080 52828 3108
rect 1544 3068 1550 3080
rect 1397 3043 1455 3049
rect 1397 3009 1409 3043
rect 1443 3040 1455 3043
rect 2222 3040 2228 3052
rect 1443 3012 2228 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 16546 3040 16574 3080
rect 5316 3012 16574 3040
rect 5316 3000 5322 3012
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 21968 3012 22201 3040
rect 21968 3000 21974 3012
rect 22189 3009 22201 3012
rect 22235 3009 22247 3043
rect 28442 3040 28448 3052
rect 28403 3012 28448 3040
rect 22189 3003 22247 3009
rect 28442 3000 28448 3012
rect 28500 3000 28506 3052
rect 30834 3000 30840 3052
rect 30892 3040 30898 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 30892 3012 32321 3040
rect 30892 3000 30898 3012
rect 32309 3009 32321 3012
rect 32355 3040 32367 3043
rect 33042 3040 33048 3052
rect 32355 3012 33048 3040
rect 32355 3009 32367 3012
rect 32309 3003 32367 3009
rect 33042 3000 33048 3012
rect 33100 3000 33106 3052
rect 34698 3000 34704 3052
rect 34756 3040 34762 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34756 3012 34989 3040
rect 34756 3000 34762 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 40037 3043 40095 3049
rect 34977 3003 35035 3009
rect 35084 3012 35572 3040
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8352 2944 8401 2972
rect 8352 2932 8358 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 32122 2972 32128 2984
rect 8389 2935 8447 2941
rect 16546 2944 26234 2972
rect 32083 2944 32128 2972
rect 1854 2864 1860 2916
rect 1912 2904 1918 2916
rect 16546 2904 16574 2944
rect 1912 2876 16574 2904
rect 26206 2904 26234 2944
rect 32122 2932 32128 2944
rect 32180 2932 32186 2984
rect 35084 2972 35112 3012
rect 34716 2944 35112 2972
rect 34716 2904 34744 2944
rect 26206 2876 34744 2904
rect 35544 2904 35572 3012
rect 40037 3009 40049 3043
rect 40083 3040 40095 3043
rect 40126 3040 40132 3052
rect 40083 3012 40132 3040
rect 40083 3009 40095 3012
rect 40037 3003 40095 3009
rect 40126 3000 40132 3012
rect 40184 3000 40190 3052
rect 43346 3040 43352 3052
rect 43307 3012 43352 3040
rect 43346 3000 43352 3012
rect 43404 3000 43410 3052
rect 43456 3040 43484 3080
rect 52822 3068 52828 3080
rect 52880 3068 52886 3120
rect 46382 3040 46388 3052
rect 43456 3012 46388 3040
rect 46382 3000 46388 3012
rect 46440 3000 46446 3052
rect 47762 3040 47768 3052
rect 47723 3012 47768 3040
rect 47762 3000 47768 3012
rect 47820 3000 47826 3052
rect 50249 3043 50307 3049
rect 50249 3040 50261 3043
rect 47872 3012 50261 3040
rect 35618 2932 35624 2984
rect 35676 2972 35682 2984
rect 39666 2972 39672 2984
rect 35676 2944 39672 2972
rect 35676 2932 35682 2944
rect 39666 2932 39672 2944
rect 39724 2932 39730 2984
rect 39850 2932 39856 2984
rect 39908 2972 39914 2984
rect 43162 2972 43168 2984
rect 39908 2944 39953 2972
rect 43123 2944 43168 2972
rect 39908 2932 39914 2944
rect 43162 2932 43168 2944
rect 43220 2932 43226 2984
rect 43622 2932 43628 2984
rect 43680 2972 43686 2984
rect 44177 2975 44235 2981
rect 44177 2972 44189 2975
rect 43680 2944 44189 2972
rect 43680 2932 43686 2944
rect 44177 2941 44189 2944
rect 44223 2941 44235 2975
rect 47578 2972 47584 2984
rect 47539 2944 47584 2972
rect 44177 2935 44235 2941
rect 47578 2932 47584 2944
rect 47636 2932 47642 2984
rect 43533 2907 43591 2913
rect 35544 2876 41414 2904
rect 1912 2864 1918 2876
rect 1118 2796 1124 2848
rect 1176 2836 1182 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1176 2808 1593 2836
rect 1176 2796 1182 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2832 2808 3065 2836
rect 2832 2796 2838 2808
rect 3053 2805 3065 2808
rect 3099 2805 3111 2839
rect 22002 2836 22008 2848
rect 21963 2808 22008 2836
rect 3053 2799 3111 2805
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 28350 2796 28356 2848
rect 28408 2836 28414 2848
rect 28629 2839 28687 2845
rect 28629 2836 28641 2839
rect 28408 2808 28641 2836
rect 28408 2796 28414 2808
rect 28629 2805 28641 2808
rect 28675 2805 28687 2839
rect 28629 2799 28687 2805
rect 29086 2796 29092 2848
rect 29144 2836 29150 2848
rect 29365 2839 29423 2845
rect 29365 2836 29377 2839
rect 29144 2808 29377 2836
rect 29144 2796 29150 2808
rect 29365 2805 29377 2808
rect 29411 2805 29423 2839
rect 31570 2836 31576 2848
rect 31531 2808 31576 2836
rect 29365 2799 29423 2805
rect 31570 2796 31576 2808
rect 31628 2796 31634 2848
rect 32493 2839 32551 2845
rect 32493 2805 32505 2839
rect 32539 2836 32551 2839
rect 32858 2836 32864 2848
rect 32539 2808 32864 2836
rect 32539 2805 32551 2808
rect 32493 2799 32551 2805
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 34793 2839 34851 2845
rect 34793 2805 34805 2839
rect 34839 2836 34851 2839
rect 35434 2836 35440 2848
rect 34839 2808 35440 2836
rect 34839 2805 34851 2808
rect 34793 2799 34851 2805
rect 35434 2796 35440 2808
rect 35492 2796 35498 2848
rect 35526 2796 35532 2848
rect 35584 2836 35590 2848
rect 35805 2839 35863 2845
rect 35805 2836 35817 2839
rect 35584 2808 35817 2836
rect 35584 2796 35590 2808
rect 35805 2805 35817 2808
rect 35851 2805 35863 2839
rect 35805 2799 35863 2805
rect 37090 2796 37096 2848
rect 37148 2836 37154 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 37148 2808 37473 2836
rect 37148 2796 37154 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 39482 2796 39488 2848
rect 39540 2836 39546 2848
rect 39761 2839 39819 2845
rect 39761 2836 39773 2839
rect 39540 2808 39773 2836
rect 39540 2796 39546 2808
rect 39761 2805 39773 2808
rect 39807 2805 39819 2839
rect 40218 2836 40224 2848
rect 40179 2808 40224 2836
rect 39761 2799 39819 2805
rect 40218 2796 40224 2808
rect 40276 2796 40282 2848
rect 41386 2836 41414 2876
rect 43533 2873 43545 2907
rect 43579 2904 43591 2907
rect 47872 2904 47900 3012
rect 50249 3009 50261 3012
rect 50295 3009 50307 3043
rect 50614 3040 50620 3052
rect 50575 3012 50620 3040
rect 50249 3003 50307 3009
rect 50614 3000 50620 3012
rect 50672 3000 50678 3052
rect 52181 3043 52239 3049
rect 52181 3009 52193 3043
rect 52227 3040 52239 3043
rect 52362 3040 52368 3052
rect 52227 3012 52368 3040
rect 52227 3009 52239 3012
rect 52181 3003 52239 3009
rect 52362 3000 52368 3012
rect 52420 3000 52426 3052
rect 52932 3049 52960 3148
rect 53282 3136 53288 3148
rect 53340 3136 53346 3188
rect 54938 3176 54944 3188
rect 54899 3148 54944 3176
rect 54938 3136 54944 3148
rect 54996 3136 55002 3188
rect 57885 3179 57943 3185
rect 57885 3176 57897 3179
rect 56704 3148 57897 3176
rect 53116 3080 55996 3108
rect 52917 3043 52975 3049
rect 52917 3009 52929 3043
rect 52963 3009 52975 3043
rect 52917 3003 52975 3009
rect 53006 3000 53012 3052
rect 53064 3040 53070 3052
rect 53116 3049 53144 3080
rect 55968 3049 55996 3080
rect 53101 3043 53159 3049
rect 53101 3040 53113 3043
rect 53064 3012 53113 3040
rect 53064 3000 53070 3012
rect 53101 3009 53113 3012
rect 53147 3009 53159 3043
rect 53101 3003 53159 3009
rect 54757 3043 54815 3049
rect 54757 3009 54769 3043
rect 54803 3009 54815 3043
rect 54757 3003 54815 3009
rect 55953 3043 56011 3049
rect 55953 3009 55965 3043
rect 55999 3040 56011 3043
rect 56594 3040 56600 3052
rect 55999 3012 56600 3040
rect 55999 3009 56011 3012
rect 55953 3003 56011 3009
rect 47949 2975 48007 2981
rect 47949 2941 47961 2975
rect 47995 2972 48007 2975
rect 54772 2972 54800 3003
rect 56594 3000 56600 3012
rect 56652 3000 56658 3052
rect 56704 3049 56732 3148
rect 57885 3145 57897 3148
rect 57931 3145 57943 3179
rect 57885 3139 57943 3145
rect 57974 3136 57980 3188
rect 58032 3176 58038 3188
rect 62390 3176 62396 3188
rect 58032 3148 62396 3176
rect 58032 3136 58038 3148
rect 62390 3136 62396 3148
rect 62448 3136 62454 3188
rect 66346 3176 66352 3188
rect 66307 3148 66352 3176
rect 66346 3136 66352 3148
rect 66404 3136 66410 3188
rect 68370 3176 68376 3188
rect 68331 3148 68376 3176
rect 68370 3136 68376 3148
rect 68428 3136 68434 3188
rect 83550 3136 83556 3188
rect 83608 3176 83614 3188
rect 112622 3176 112628 3188
rect 83608 3148 112628 3176
rect 83608 3136 83614 3148
rect 112622 3136 112628 3148
rect 112680 3136 112686 3188
rect 113361 3179 113419 3185
rect 113361 3176 113373 3179
rect 113146 3148 113373 3176
rect 56962 3108 56968 3120
rect 56923 3080 56968 3108
rect 56962 3068 56968 3080
rect 57020 3068 57026 3120
rect 61838 3068 61844 3120
rect 61896 3108 61902 3120
rect 61896 3080 63264 3108
rect 61896 3068 61902 3080
rect 56689 3043 56747 3049
rect 56689 3009 56701 3043
rect 56735 3009 56747 3043
rect 56689 3003 56747 3009
rect 56778 3000 56784 3052
rect 56836 3040 56842 3052
rect 56836 3012 56881 3040
rect 56836 3000 56842 3012
rect 57146 3000 57152 3052
rect 57204 3040 57210 3052
rect 58069 3043 58127 3049
rect 58069 3040 58081 3043
rect 57204 3012 58081 3040
rect 57204 3000 57210 3012
rect 58069 3009 58081 3012
rect 58115 3009 58127 3043
rect 58069 3003 58127 3009
rect 59538 3000 59544 3052
rect 59596 3040 59602 3052
rect 59817 3043 59875 3049
rect 59817 3040 59829 3043
rect 59596 3012 59829 3040
rect 59596 3000 59602 3012
rect 59817 3009 59829 3012
rect 59863 3009 59875 3043
rect 59817 3003 59875 3009
rect 61105 3043 61163 3049
rect 61105 3009 61117 3043
rect 61151 3040 61163 3043
rect 61930 3040 61936 3052
rect 61151 3012 61936 3040
rect 61151 3009 61163 3012
rect 61105 3003 61163 3009
rect 61930 3000 61936 3012
rect 61988 3000 61994 3052
rect 63236 3049 63264 3080
rect 79134 3068 79140 3120
rect 79192 3108 79198 3120
rect 83921 3111 83979 3117
rect 83921 3108 83933 3111
rect 79192 3080 83933 3108
rect 79192 3068 79198 3080
rect 83921 3077 83933 3080
rect 83967 3077 83979 3111
rect 83921 3071 83979 3077
rect 84856 3080 89300 3108
rect 63221 3043 63279 3049
rect 63221 3009 63233 3043
rect 63267 3009 63279 3043
rect 66254 3040 66260 3052
rect 66215 3012 66260 3040
rect 63221 3003 63279 3009
rect 66254 3000 66260 3012
rect 66312 3000 66318 3052
rect 68186 3040 68192 3052
rect 68147 3012 68192 3040
rect 68186 3000 68192 3012
rect 68244 3000 68250 3052
rect 69293 3043 69351 3049
rect 69293 3009 69305 3043
rect 69339 3040 69351 3043
rect 70581 3043 70639 3049
rect 70581 3040 70593 3043
rect 69339 3012 70593 3040
rect 69339 3009 69351 3012
rect 69293 3003 69351 3009
rect 70581 3009 70593 3012
rect 70627 3040 70639 3043
rect 73614 3040 73620 3052
rect 70627 3012 71452 3040
rect 73575 3012 73620 3040
rect 70627 3009 70639 3012
rect 70581 3003 70639 3009
rect 47995 2944 54800 2972
rect 47995 2941 48007 2944
rect 47949 2935 48007 2941
rect 54846 2932 54852 2984
rect 54904 2972 54910 2984
rect 55769 2975 55827 2981
rect 55769 2972 55781 2975
rect 54904 2944 55781 2972
rect 54904 2932 54910 2944
rect 55769 2941 55781 2944
rect 55815 2941 55827 2975
rect 55769 2935 55827 2941
rect 56137 2975 56195 2981
rect 56137 2941 56149 2975
rect 56183 2972 56195 2975
rect 57330 2972 57336 2984
rect 56183 2944 57336 2972
rect 56183 2941 56195 2944
rect 56137 2935 56195 2941
rect 57330 2932 57336 2944
rect 57388 2932 57394 2984
rect 61841 2975 61899 2981
rect 61841 2972 61853 2975
rect 57532 2944 61853 2972
rect 57422 2904 57428 2916
rect 43579 2876 47900 2904
rect 47964 2876 57428 2904
rect 43579 2873 43591 2876
rect 43533 2867 43591 2873
rect 46198 2836 46204 2848
rect 41386 2808 46204 2836
rect 46198 2796 46204 2808
rect 46256 2796 46262 2848
rect 46290 2796 46296 2848
rect 46348 2836 46354 2848
rect 47964 2836 47992 2876
rect 57422 2864 57428 2876
rect 57480 2864 57486 2916
rect 46348 2808 47992 2836
rect 46348 2796 46354 2808
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51261 2839 51319 2845
rect 51261 2836 51273 2839
rect 50764 2808 51273 2836
rect 50764 2796 50770 2808
rect 51261 2805 51273 2808
rect 51307 2805 51319 2839
rect 51261 2799 51319 2805
rect 51902 2796 51908 2848
rect 51960 2836 51966 2848
rect 57532 2836 57560 2944
rect 61841 2941 61853 2944
rect 61887 2941 61899 2975
rect 61841 2935 61899 2941
rect 68646 2932 68652 2984
rect 68704 2972 68710 2984
rect 69569 2975 69627 2981
rect 69569 2972 69581 2975
rect 68704 2944 69581 2972
rect 68704 2932 68710 2944
rect 69569 2941 69581 2944
rect 69615 2941 69627 2975
rect 70762 2972 70768 2984
rect 70723 2944 70768 2972
rect 69569 2935 69627 2941
rect 70762 2932 70768 2944
rect 70820 2932 70826 2984
rect 71424 2972 71452 3012
rect 73614 3000 73620 3012
rect 73672 3000 73678 3052
rect 73706 3000 73712 3052
rect 73764 3040 73770 3052
rect 74353 3043 74411 3049
rect 74353 3040 74365 3043
rect 73764 3012 74365 3040
rect 73764 3000 73770 3012
rect 74353 3009 74365 3012
rect 74399 3009 74411 3043
rect 74353 3003 74411 3009
rect 76282 3000 76288 3052
rect 76340 3040 76346 3052
rect 76561 3043 76619 3049
rect 76561 3040 76573 3043
rect 76340 3012 76573 3040
rect 76340 3000 76346 3012
rect 76561 3009 76573 3012
rect 76607 3009 76619 3043
rect 76561 3003 76619 3009
rect 76742 3000 76748 3052
rect 76800 3040 76806 3052
rect 79689 3043 79747 3049
rect 79689 3040 79701 3043
rect 76800 3012 79701 3040
rect 76800 3000 76806 3012
rect 79689 3009 79701 3012
rect 79735 3040 79747 3043
rect 83642 3040 83648 3052
rect 79735 3012 83504 3040
rect 83603 3012 83648 3040
rect 79735 3009 79747 3012
rect 79689 3003 79747 3009
rect 76760 2972 76788 3000
rect 79962 2972 79968 2984
rect 71424 2944 76788 2972
rect 79923 2944 79968 2972
rect 79962 2932 79968 2944
rect 80020 2932 80026 2984
rect 83476 2972 83504 3012
rect 83642 3000 83648 3012
rect 83700 3000 83706 3052
rect 84856 2972 84884 3080
rect 85942 3000 85948 3052
rect 86000 3040 86006 3052
rect 86221 3043 86279 3049
rect 86221 3040 86233 3043
rect 86000 3012 86233 3040
rect 86000 3000 86006 3012
rect 86221 3009 86233 3012
rect 86267 3009 86279 3043
rect 86221 3003 86279 3009
rect 86589 3043 86647 3049
rect 86589 3009 86601 3043
rect 86635 3040 86647 3043
rect 86862 3040 86868 3052
rect 86635 3012 86868 3040
rect 86635 3009 86647 3012
rect 86589 3003 86647 3009
rect 86862 3000 86868 3012
rect 86920 3000 86926 3052
rect 87417 3043 87475 3049
rect 87417 3009 87429 3043
rect 87463 3040 87475 3043
rect 88150 3040 88156 3052
rect 87463 3012 88156 3040
rect 87463 3009 87475 3012
rect 87417 3003 87475 3009
rect 88150 3000 88156 3012
rect 88208 3000 88214 3052
rect 83476 2944 84884 2972
rect 86880 2972 86908 3000
rect 87601 2975 87659 2981
rect 87601 2972 87613 2975
rect 86880 2944 87613 2972
rect 87601 2941 87613 2944
rect 87647 2972 87659 2975
rect 88981 2975 89039 2981
rect 88981 2972 88993 2975
rect 87647 2944 88993 2972
rect 87647 2941 87659 2944
rect 87601 2935 87659 2941
rect 88981 2941 88993 2944
rect 89027 2941 89039 2975
rect 88981 2935 89039 2941
rect 89165 2975 89223 2981
rect 89165 2941 89177 2975
rect 89211 2941 89223 2975
rect 89272 2972 89300 3080
rect 89622 3068 89628 3120
rect 89680 3108 89686 3120
rect 93854 3108 93860 3120
rect 89680 3080 93860 3108
rect 89680 3068 89686 3080
rect 93854 3068 93860 3080
rect 93912 3068 93918 3120
rect 94216 3111 94274 3117
rect 94216 3077 94228 3111
rect 94262 3108 94274 3111
rect 94958 3108 94964 3120
rect 94262 3080 94964 3108
rect 94262 3077 94274 3080
rect 94216 3071 94274 3077
rect 94958 3068 94964 3080
rect 95016 3068 95022 3120
rect 95050 3068 95056 3120
rect 95108 3108 95114 3120
rect 100849 3111 100907 3117
rect 95108 3080 100432 3108
rect 95108 3068 95114 3080
rect 100404 3052 100432 3080
rect 100849 3077 100861 3111
rect 100895 3108 100907 3111
rect 111788 3111 111846 3117
rect 100895 3080 110920 3108
rect 100895 3077 100907 3080
rect 100849 3071 100907 3077
rect 89346 3000 89352 3052
rect 89404 3040 89410 3052
rect 89533 3043 89591 3049
rect 89404 3012 89449 3040
rect 89404 3000 89410 3012
rect 89533 3009 89545 3043
rect 89579 3040 89591 3043
rect 90177 3043 90235 3049
rect 90177 3040 90189 3043
rect 89579 3012 90189 3040
rect 89579 3009 89591 3012
rect 89533 3003 89591 3009
rect 90177 3009 90189 3012
rect 90223 3009 90235 3043
rect 91186 3040 91192 3052
rect 91147 3012 91192 3040
rect 90177 3003 90235 3009
rect 91186 3000 91192 3012
rect 91244 3000 91250 3052
rect 92014 3040 92020 3052
rect 91975 3012 92020 3040
rect 92014 3000 92020 3012
rect 92072 3000 92078 3052
rect 93949 3043 94007 3049
rect 93949 3009 93961 3043
rect 93995 3040 94007 3043
rect 94038 3040 94044 3052
rect 93995 3012 94044 3040
rect 93995 3009 94007 3012
rect 93949 3003 94007 3009
rect 94038 3000 94044 3012
rect 94096 3000 94102 3052
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 97077 3043 97135 3049
rect 97077 3040 97089 3043
rect 96948 3012 97089 3040
rect 96948 3000 96954 3012
rect 97077 3009 97089 3012
rect 97123 3009 97135 3043
rect 99558 3040 99564 3052
rect 99471 3012 99564 3040
rect 97077 3003 97135 3009
rect 99558 3000 99564 3012
rect 99616 3040 99622 3052
rect 100113 3043 100171 3049
rect 100113 3040 100125 3043
rect 99616 3012 100125 3040
rect 99616 3000 99622 3012
rect 100113 3009 100125 3012
rect 100159 3009 100171 3043
rect 100113 3003 100171 3009
rect 100386 3000 100392 3052
rect 100444 3040 100450 3052
rect 100757 3043 100815 3049
rect 100757 3040 100769 3043
rect 100444 3012 100769 3040
rect 100444 3000 100450 3012
rect 100757 3009 100769 3012
rect 100803 3009 100815 3043
rect 104250 3040 104256 3052
rect 104211 3012 104256 3040
rect 100757 3003 100815 3009
rect 104250 3000 104256 3012
rect 104308 3000 104314 3052
rect 104986 3000 104992 3052
rect 105044 3040 105050 3052
rect 105173 3043 105231 3049
rect 105173 3040 105185 3043
rect 105044 3012 105185 3040
rect 105044 3000 105050 3012
rect 105173 3009 105185 3012
rect 105219 3009 105231 3043
rect 107286 3040 107292 3052
rect 107247 3012 107292 3040
rect 105173 3003 105231 3009
rect 107286 3000 107292 3012
rect 107344 3000 107350 3052
rect 107556 3043 107614 3049
rect 107556 3009 107568 3043
rect 107602 3040 107614 3043
rect 108298 3040 108304 3052
rect 107602 3012 108304 3040
rect 107602 3009 107614 3012
rect 107556 3003 107614 3009
rect 108298 3000 108304 3012
rect 108356 3000 108362 3052
rect 91204 2972 91232 3000
rect 89272 2944 91232 2972
rect 89165 2935 89223 2941
rect 57606 2864 57612 2916
rect 57664 2904 57670 2916
rect 73801 2907 73859 2913
rect 73801 2904 73813 2907
rect 57664 2876 73813 2904
rect 57664 2864 57670 2876
rect 73801 2873 73813 2876
rect 73847 2873 73859 2907
rect 73801 2867 73859 2873
rect 73982 2864 73988 2916
rect 74040 2904 74046 2916
rect 86037 2907 86095 2913
rect 74040 2876 84516 2904
rect 74040 2864 74046 2876
rect 51960 2808 57560 2836
rect 59633 2839 59691 2845
rect 51960 2796 51966 2808
rect 59633 2805 59645 2839
rect 59679 2836 59691 2839
rect 62022 2836 62028 2848
rect 59679 2808 62028 2836
rect 59679 2805 59691 2808
rect 59633 2799 59691 2805
rect 62022 2796 62028 2808
rect 62080 2796 62086 2848
rect 62114 2796 62120 2848
rect 62172 2836 62178 2848
rect 63037 2839 63095 2845
rect 63037 2836 63049 2839
rect 62172 2808 63049 2836
rect 62172 2796 62178 2808
rect 63037 2805 63049 2808
rect 63083 2805 63095 2839
rect 63037 2799 63095 2805
rect 65150 2796 65156 2848
rect 65208 2836 65214 2848
rect 65429 2839 65487 2845
rect 65429 2836 65441 2839
rect 65208 2808 65441 2836
rect 65208 2796 65214 2808
rect 65429 2805 65441 2808
rect 65475 2805 65487 2839
rect 65429 2799 65487 2805
rect 74537 2839 74595 2845
rect 74537 2805 74549 2839
rect 74583 2836 74595 2839
rect 74626 2836 74632 2848
rect 74583 2808 74632 2836
rect 74583 2805 74595 2808
rect 74537 2799 74595 2805
rect 74626 2796 74632 2808
rect 74684 2796 74690 2848
rect 74718 2796 74724 2848
rect 74776 2836 74782 2848
rect 75273 2839 75331 2845
rect 75273 2836 75285 2839
rect 74776 2808 75285 2836
rect 74776 2796 74782 2808
rect 75273 2805 75285 2808
rect 75319 2805 75331 2839
rect 76374 2836 76380 2848
rect 76335 2808 76380 2836
rect 75273 2799 75331 2805
rect 76374 2796 76380 2808
rect 76432 2796 76438 2848
rect 77110 2796 77116 2848
rect 77168 2836 77174 2848
rect 77389 2839 77447 2845
rect 77389 2836 77401 2839
rect 77168 2808 77401 2836
rect 77168 2796 77174 2808
rect 77389 2805 77401 2808
rect 77435 2805 77447 2839
rect 77389 2799 77447 2805
rect 81894 2796 81900 2848
rect 81952 2836 81958 2848
rect 82173 2839 82231 2845
rect 82173 2836 82185 2839
rect 81952 2808 82185 2836
rect 81952 2796 81958 2808
rect 82173 2805 82185 2808
rect 82219 2805 82231 2839
rect 84488 2836 84516 2876
rect 86037 2873 86049 2907
rect 86083 2904 86095 2907
rect 89180 2904 89208 2935
rect 97994 2932 98000 2984
rect 98052 2972 98058 2984
rect 101033 2975 101091 2981
rect 101033 2972 101045 2975
rect 98052 2944 101045 2972
rect 98052 2932 98058 2944
rect 101033 2941 101045 2944
rect 101079 2972 101091 2975
rect 101079 2944 105492 2972
rect 101079 2941 101091 2944
rect 101033 2935 101091 2941
rect 90634 2904 90640 2916
rect 86083 2876 89208 2904
rect 89364 2876 90640 2904
rect 86083 2873 86095 2876
rect 86037 2867 86095 2873
rect 89364 2848 89392 2876
rect 90634 2864 90640 2876
rect 90692 2904 90698 2916
rect 91005 2907 91063 2913
rect 91005 2904 91017 2907
rect 90692 2876 91017 2904
rect 90692 2864 90698 2876
rect 91005 2873 91017 2876
rect 91051 2873 91063 2907
rect 91005 2867 91063 2873
rect 91738 2864 91744 2916
rect 91796 2904 91802 2916
rect 96982 2904 96988 2916
rect 91796 2876 93992 2904
rect 91796 2864 91802 2876
rect 87690 2836 87696 2848
rect 84488 2808 87696 2836
rect 82173 2799 82231 2805
rect 87690 2796 87696 2808
rect 87748 2796 87754 2848
rect 87966 2796 87972 2848
rect 88024 2836 88030 2848
rect 89346 2836 89352 2848
rect 88024 2808 89352 2836
rect 88024 2796 88030 2808
rect 89346 2796 89352 2808
rect 89404 2796 89410 2848
rect 90266 2836 90272 2848
rect 90227 2808 90272 2836
rect 90266 2796 90272 2808
rect 90324 2796 90330 2848
rect 92106 2836 92112 2848
rect 92067 2808 92112 2836
rect 92106 2796 92112 2808
rect 92164 2796 92170 2848
rect 93964 2836 93992 2876
rect 95344 2876 96988 2904
rect 95344 2845 95372 2876
rect 96982 2864 96988 2876
rect 97040 2864 97046 2916
rect 97261 2907 97319 2913
rect 97261 2873 97273 2907
rect 97307 2904 97319 2907
rect 105170 2904 105176 2916
rect 97307 2876 105176 2904
rect 97307 2873 97319 2876
rect 97261 2867 97319 2873
rect 105170 2864 105176 2876
rect 105228 2864 105234 2916
rect 95329 2839 95387 2845
rect 95329 2836 95341 2839
rect 93964 2808 95341 2836
rect 95329 2805 95341 2808
rect 95375 2805 95387 2839
rect 95329 2799 95387 2805
rect 96246 2796 96252 2848
rect 96304 2836 96310 2848
rect 96617 2839 96675 2845
rect 96617 2836 96629 2839
rect 96304 2808 96629 2836
rect 96304 2796 96310 2808
rect 96617 2805 96629 2808
rect 96663 2805 96675 2839
rect 96617 2799 96675 2805
rect 99466 2796 99472 2848
rect 99524 2836 99530 2848
rect 99745 2839 99803 2845
rect 99745 2836 99757 2839
rect 99524 2808 99757 2836
rect 99524 2796 99530 2808
rect 99745 2805 99757 2808
rect 99791 2805 99803 2839
rect 99745 2799 99803 2805
rect 100389 2839 100447 2845
rect 100389 2805 100401 2839
rect 100435 2836 100447 2839
rect 100938 2836 100944 2848
rect 100435 2808 100944 2836
rect 100435 2805 100447 2808
rect 100389 2799 100447 2805
rect 100938 2796 100944 2808
rect 100996 2796 101002 2848
rect 103514 2796 103520 2848
rect 103572 2836 103578 2848
rect 104437 2839 104495 2845
rect 104437 2836 104449 2839
rect 103572 2808 104449 2836
rect 103572 2796 103578 2808
rect 104437 2805 104449 2808
rect 104483 2805 104495 2839
rect 104437 2799 104495 2805
rect 105078 2796 105084 2848
rect 105136 2836 105142 2848
rect 105357 2839 105415 2845
rect 105357 2836 105369 2839
rect 105136 2808 105369 2836
rect 105136 2796 105142 2808
rect 105357 2805 105369 2808
rect 105403 2805 105415 2839
rect 105464 2836 105492 2944
rect 108669 2907 108727 2913
rect 108669 2873 108681 2907
rect 108715 2904 108727 2907
rect 109770 2904 109776 2916
rect 108715 2876 109776 2904
rect 108715 2873 108727 2876
rect 108669 2867 108727 2873
rect 109770 2864 109776 2876
rect 109828 2864 109834 2916
rect 110892 2913 110920 3080
rect 111788 3077 111800 3111
rect 111834 3108 111846 3111
rect 113146 3108 113174 3148
rect 113361 3145 113373 3148
rect 113407 3145 113419 3179
rect 113361 3139 113419 3145
rect 115566 3136 115572 3188
rect 115624 3176 115630 3188
rect 118053 3179 118111 3185
rect 118053 3176 118065 3179
rect 115624 3148 118065 3176
rect 115624 3136 115630 3148
rect 118053 3145 118065 3148
rect 118099 3145 118111 3179
rect 118053 3139 118111 3145
rect 111834 3080 113174 3108
rect 111834 3077 111846 3080
rect 111788 3071 111846 3077
rect 111061 3043 111119 3049
rect 111061 3009 111073 3043
rect 111107 3040 111119 3043
rect 111426 3040 111432 3052
rect 111107 3012 111432 3040
rect 111107 3009 111119 3012
rect 111061 3003 111119 3009
rect 111426 3000 111432 3012
rect 111484 3000 111490 3052
rect 112254 3000 112260 3052
rect 112312 3040 112318 3052
rect 113545 3043 113603 3049
rect 113545 3040 113557 3043
rect 112312 3012 113557 3040
rect 112312 3000 112318 3012
rect 113545 3009 113557 3012
rect 113591 3009 113603 3043
rect 114830 3040 114836 3052
rect 114791 3012 114836 3040
rect 113545 3003 113603 3009
rect 114830 3000 114836 3012
rect 114888 3000 114894 3052
rect 117958 3040 117964 3052
rect 117919 3012 117964 3040
rect 117958 3000 117964 3012
rect 118016 3000 118022 3052
rect 110966 2932 110972 2984
rect 111024 2972 111030 2984
rect 111521 2975 111579 2981
rect 111521 2972 111533 2975
rect 111024 2944 111533 2972
rect 111024 2932 111030 2944
rect 111521 2941 111533 2944
rect 111567 2941 111579 2975
rect 111521 2935 111579 2941
rect 110877 2907 110935 2913
rect 110877 2873 110889 2907
rect 110923 2873 110935 2907
rect 110877 2867 110935 2873
rect 109954 2836 109960 2848
rect 105464 2808 109960 2836
rect 105357 2799 105415 2805
rect 109954 2796 109960 2808
rect 110012 2796 110018 2848
rect 112162 2796 112168 2848
rect 112220 2836 112226 2848
rect 112901 2839 112959 2845
rect 112901 2836 112913 2839
rect 112220 2808 112913 2836
rect 112220 2796 112226 2808
rect 112901 2805 112913 2808
rect 112947 2805 112959 2839
rect 112901 2799 112959 2805
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 115017 2839 115075 2845
rect 115017 2836 115029 2839
rect 114796 2808 115029 2836
rect 114796 2796 114802 2808
rect 115017 2805 115029 2808
rect 115063 2805 115075 2839
rect 115017 2799 115075 2805
rect 1104 2746 118864 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 118864 2746
rect 1104 2672 118864 2694
rect 22370 2632 22376 2644
rect 22331 2604 22376 2632
rect 22370 2592 22376 2604
rect 22428 2592 22434 2644
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 28626 2632 28632 2644
rect 23532 2604 28632 2632
rect 23532 2592 23538 2604
rect 28626 2592 28632 2604
rect 28684 2632 28690 2644
rect 30834 2632 30840 2644
rect 28684 2604 30840 2632
rect 28684 2592 28690 2604
rect 30834 2592 30840 2604
rect 30892 2592 30898 2644
rect 37826 2632 37832 2644
rect 30944 2604 37832 2632
rect 30944 2564 30972 2604
rect 37826 2592 37832 2604
rect 37884 2592 37890 2644
rect 43162 2632 43168 2644
rect 39500 2604 43168 2632
rect 14844 2536 30972 2564
rect 2406 2496 2412 2508
rect 2367 2468 2412 2496
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 4338 2388 4344 2440
rect 4396 2428 4402 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4396 2400 4629 2428
rect 4396 2388 4402 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5258 2428 5264 2440
rect 5031 2400 5264 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5902 2388 5908 2440
rect 5960 2428 5966 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5960 2400 6561 2428
rect 5960 2388 5966 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 9180 2400 9413 2428
rect 9180 2388 9186 2400
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 9401 2391 9459 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10778 2388 10784 2440
rect 10836 2428 10842 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 10836 2400 11713 2428
rect 10836 2388 10842 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 13906 2428 13912 2440
rect 13867 2400 13912 2428
rect 11701 2391 11759 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 14844 2437 14872 2536
rect 33134 2524 33140 2576
rect 33192 2564 33198 2576
rect 33965 2567 34023 2573
rect 33965 2564 33977 2567
rect 33192 2536 33977 2564
rect 33192 2524 33198 2536
rect 33965 2533 33977 2536
rect 34011 2533 34023 2567
rect 39500 2564 39528 2604
rect 43162 2592 43168 2604
rect 43220 2592 43226 2644
rect 43254 2592 43260 2644
rect 43312 2632 43318 2644
rect 43717 2635 43775 2641
rect 43312 2604 43484 2632
rect 43312 2592 43318 2604
rect 33965 2527 34023 2533
rect 34164 2536 39528 2564
rect 42705 2567 42763 2573
rect 34054 2496 34060 2508
rect 16546 2468 34060 2496
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14599 2400 14841 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15620 2400 15853 2428
rect 15620 2388 15626 2400
rect 15841 2397 15853 2400
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 7745 2363 7803 2369
rect 7745 2360 7757 2363
rect 7616 2332 7757 2360
rect 7616 2320 7622 2332
rect 7745 2329 7757 2332
rect 7791 2329 7803 2363
rect 7745 2323 7803 2329
rect 12342 2320 12348 2372
rect 12400 2360 12406 2372
rect 12529 2363 12587 2369
rect 12529 2360 12541 2363
rect 12400 2332 12541 2360
rect 12400 2320 12406 2332
rect 12529 2329 12541 2332
rect 12575 2329 12587 2363
rect 12529 2323 12587 2329
rect 12713 2363 12771 2369
rect 12713 2329 12725 2363
rect 12759 2360 12771 2363
rect 16546 2360 16574 2468
rect 34054 2456 34060 2468
rect 34112 2456 34118 2508
rect 17126 2388 17132 2440
rect 17184 2428 17190 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 17184 2400 17417 2428
rect 17184 2388 17190 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 18690 2428 18696 2440
rect 18651 2400 18696 2428
rect 17405 2391 17463 2397
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 19426 2388 19432 2440
rect 19484 2428 19490 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19484 2400 19625 2428
rect 19484 2388 19490 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20404 2400 20637 2428
rect 20404 2388 20410 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 22002 2428 22008 2440
rect 21963 2400 22008 2428
rect 20625 2391 20683 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 23474 2428 23480 2440
rect 22235 2400 23480 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23624 2400 23857 2428
rect 23624 2388 23630 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 24394 2428 24400 2440
rect 24355 2400 24400 2428
rect 23845 2391 23903 2397
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25409 2431 25467 2437
rect 25409 2428 25421 2431
rect 25188 2400 25421 2428
rect 25188 2388 25194 2400
rect 25409 2397 25421 2400
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 26694 2388 26700 2440
rect 26752 2428 26758 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26752 2400 27169 2428
rect 26752 2388 26758 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27522 2388 27528 2440
rect 27580 2428 27586 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27580 2400 27813 2428
rect 27580 2388 27586 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28445 2431 28503 2437
rect 28445 2397 28457 2431
rect 28491 2397 28503 2431
rect 28626 2428 28632 2440
rect 28587 2400 28632 2428
rect 28445 2391 28503 2397
rect 26878 2360 26884 2372
rect 12759 2332 16574 2360
rect 17236 2332 26884 2360
rect 12759 2329 12771 2332
rect 12713 2323 12771 2329
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3568 2264 3801 2292
rect 3568 2252 3574 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 7834 2292 7840 2304
rect 7795 2264 7840 2292
rect 5445 2255 5503 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 9950 2252 9956 2304
rect 10008 2292 10014 2304
rect 10229 2295 10287 2301
rect 10229 2292 10241 2295
rect 10008 2264 10241 2292
rect 10008 2252 10014 2264
rect 10229 2261 10241 2264
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13228 2264 13277 2292
rect 13228 2252 13234 2264
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 17236 2301 17264 2332
rect 26878 2320 26884 2332
rect 26936 2320 26942 2372
rect 28460 2360 28488 2391
rect 28626 2388 28632 2400
rect 28684 2388 28690 2440
rect 28813 2431 28871 2437
rect 28813 2397 28825 2431
rect 28859 2428 28871 2431
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 28859 2400 29561 2428
rect 28859 2397 28871 2400
rect 28813 2391 28871 2397
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31389 2431 31447 2437
rect 31389 2397 31401 2431
rect 31435 2428 31447 2431
rect 31662 2428 31668 2440
rect 31435 2400 31668 2428
rect 31435 2397 31447 2400
rect 31389 2391 31447 2397
rect 31662 2388 31668 2400
rect 31720 2388 31726 2440
rect 32858 2428 32864 2440
rect 32819 2400 32864 2428
rect 32858 2388 32864 2400
rect 32916 2388 32922 2440
rect 34164 2428 34192 2536
rect 42705 2533 42717 2567
rect 42751 2564 42763 2567
rect 43456 2564 43484 2604
rect 43717 2601 43729 2635
rect 43763 2632 43775 2635
rect 45462 2632 45468 2644
rect 43763 2604 45468 2632
rect 43763 2601 43775 2604
rect 43717 2595 43775 2601
rect 45462 2592 45468 2604
rect 45520 2592 45526 2644
rect 49421 2635 49479 2641
rect 49421 2601 49433 2635
rect 49467 2632 49479 2635
rect 52270 2632 52276 2644
rect 49467 2604 52276 2632
rect 49467 2601 49479 2604
rect 49421 2595 49479 2601
rect 52270 2592 52276 2604
rect 52328 2592 52334 2644
rect 52454 2592 52460 2644
rect 52512 2632 52518 2644
rect 53101 2635 53159 2641
rect 53101 2632 53113 2635
rect 52512 2604 53113 2632
rect 52512 2592 52518 2604
rect 53101 2601 53113 2604
rect 53147 2601 53159 2635
rect 53101 2595 53159 2601
rect 53190 2592 53196 2644
rect 53248 2632 53254 2644
rect 85390 2632 85396 2644
rect 53248 2604 84884 2632
rect 85351 2604 85396 2632
rect 53248 2592 53254 2604
rect 61746 2564 61752 2576
rect 42751 2536 43392 2564
rect 43456 2536 61752 2564
rect 42751 2533 42763 2536
rect 42705 2527 42763 2533
rect 34238 2456 34244 2508
rect 34296 2496 34302 2508
rect 39850 2496 39856 2508
rect 34296 2468 39856 2496
rect 34296 2456 34302 2468
rect 39850 2456 39856 2468
rect 39908 2456 39914 2508
rect 43254 2496 43260 2508
rect 40236 2468 43260 2496
rect 34974 2428 34980 2440
rect 33060 2400 34192 2428
rect 34935 2400 34980 2428
rect 26988 2332 28488 2360
rect 29181 2363 29239 2369
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14792 2264 15025 2292
rect 14792 2252 14798 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2292 17923 2295
rect 17954 2292 17960 2304
rect 17911 2264 17960 2292
rect 17911 2261 17923 2264
rect 17865 2255 17923 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 19797 2295 19855 2301
rect 19797 2292 19809 2295
rect 19484 2264 19809 2292
rect 19484 2252 19490 2264
rect 19797 2261 19809 2264
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 22738 2252 22744 2304
rect 22796 2292 22802 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22796 2264 22845 2292
rect 22796 2252 22802 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 24302 2252 24308 2304
rect 24360 2292 24366 2304
rect 26988 2301 27016 2332
rect 29181 2329 29193 2363
rect 29227 2360 29239 2363
rect 29825 2363 29883 2369
rect 29825 2360 29837 2363
rect 29227 2332 29837 2360
rect 29227 2329 29239 2332
rect 29181 2323 29239 2329
rect 29825 2329 29837 2332
rect 29871 2360 29883 2363
rect 33060 2360 33088 2400
rect 34974 2388 34980 2400
rect 35032 2388 35038 2440
rect 35161 2431 35219 2437
rect 35161 2428 35173 2431
rect 35084 2400 35173 2428
rect 35084 2372 35112 2400
rect 35161 2397 35173 2400
rect 35207 2397 35219 2431
rect 35161 2391 35219 2397
rect 35345 2431 35403 2437
rect 35345 2397 35357 2431
rect 35391 2428 35403 2431
rect 36265 2431 36323 2437
rect 36265 2428 36277 2431
rect 35391 2400 36277 2428
rect 35391 2397 35403 2400
rect 35345 2391 35403 2397
rect 36265 2397 36277 2400
rect 36311 2397 36323 2431
rect 36265 2391 36323 2397
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2428 38623 2431
rect 38746 2428 38752 2440
rect 38611 2400 38752 2428
rect 38611 2397 38623 2400
rect 38565 2391 38623 2397
rect 29871 2332 30420 2360
rect 29871 2329 29883 2332
rect 29825 2323 29883 2329
rect 30392 2301 30420 2332
rect 30852 2332 33088 2360
rect 33137 2363 33195 2369
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24360 2264 24593 2292
rect 24360 2252 24366 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 26973 2295 27031 2301
rect 26973 2261 26985 2295
rect 27019 2261 27031 2295
rect 26973 2255 27031 2261
rect 30377 2295 30435 2301
rect 30377 2261 30389 2295
rect 30423 2292 30435 2295
rect 30650 2292 30656 2304
rect 30423 2264 30656 2292
rect 30423 2261 30435 2264
rect 30377 2255 30435 2261
rect 30650 2252 30656 2264
rect 30708 2252 30714 2304
rect 30852 2301 30880 2332
rect 33137 2329 33149 2363
rect 33183 2329 33195 2363
rect 33137 2323 33195 2329
rect 30837 2295 30895 2301
rect 30837 2261 30849 2295
rect 30883 2261 30895 2295
rect 30837 2255 30895 2261
rect 31849 2295 31907 2301
rect 31849 2261 31861 2295
rect 31895 2292 31907 2295
rect 32306 2292 32312 2304
rect 31895 2264 32312 2292
rect 31895 2261 31907 2264
rect 31849 2255 31907 2261
rect 32306 2252 32312 2264
rect 32364 2252 32370 2304
rect 32585 2295 32643 2301
rect 32585 2261 32597 2295
rect 32631 2292 32643 2295
rect 33152 2292 33180 2323
rect 33226 2320 33232 2372
rect 33284 2360 33290 2372
rect 35066 2360 35072 2372
rect 33284 2332 35072 2360
rect 33284 2320 33290 2332
rect 35066 2320 35072 2332
rect 35124 2320 35130 2372
rect 35989 2363 36047 2369
rect 35989 2329 36001 2363
rect 36035 2360 36047 2363
rect 36538 2360 36544 2372
rect 36035 2332 36544 2360
rect 36035 2329 36047 2332
rect 35989 2323 36047 2329
rect 36538 2320 36544 2332
rect 36596 2320 36602 2372
rect 37292 2360 37320 2391
rect 38746 2388 38752 2400
rect 38804 2388 38810 2440
rect 40236 2428 40264 2468
rect 43254 2456 43260 2468
rect 43312 2456 43318 2508
rect 43364 2505 43392 2536
rect 61746 2524 61752 2536
rect 61804 2524 61810 2576
rect 61930 2564 61936 2576
rect 61891 2536 61936 2564
rect 61930 2524 61936 2536
rect 61988 2524 61994 2576
rect 62022 2524 62028 2576
rect 62080 2564 62086 2576
rect 63405 2567 63463 2573
rect 62080 2536 63080 2564
rect 62080 2524 62086 2536
rect 43349 2499 43407 2505
rect 43349 2465 43361 2499
rect 43395 2465 43407 2499
rect 62666 2496 62672 2508
rect 43349 2459 43407 2465
rect 44376 2468 62672 2496
rect 39040 2400 40264 2428
rect 40405 2431 40463 2437
rect 37921 2363 37979 2369
rect 37921 2360 37933 2363
rect 37292 2332 37933 2360
rect 37921 2329 37933 2332
rect 37967 2360 37979 2363
rect 39040 2360 39068 2400
rect 40405 2397 40417 2431
rect 40451 2428 40463 2431
rect 40678 2428 40684 2440
rect 40451 2400 40684 2428
rect 40451 2397 40463 2400
rect 40405 2391 40463 2397
rect 40678 2388 40684 2400
rect 40736 2388 40742 2440
rect 41138 2388 41144 2440
rect 41196 2428 41202 2440
rect 41601 2431 41659 2437
rect 41601 2428 41613 2431
rect 41196 2400 41613 2428
rect 41196 2388 41202 2400
rect 41601 2397 41613 2400
rect 41647 2397 41659 2431
rect 41601 2391 41659 2397
rect 42702 2388 42708 2440
rect 42760 2428 42766 2440
rect 42889 2431 42947 2437
rect 42889 2428 42901 2431
rect 42760 2400 42901 2428
rect 42760 2388 42766 2400
rect 42889 2397 42901 2400
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 43496 2400 43545 2428
rect 43496 2388 43502 2400
rect 43533 2397 43545 2400
rect 43579 2428 43591 2431
rect 44082 2428 44088 2440
rect 43579 2400 44088 2428
rect 43579 2397 43591 2400
rect 43533 2391 43591 2397
rect 44082 2388 44088 2400
rect 44140 2388 44146 2440
rect 44376 2437 44404 2468
rect 44361 2431 44419 2437
rect 44361 2397 44373 2431
rect 44407 2397 44419 2431
rect 44361 2391 44419 2397
rect 37967 2332 39068 2360
rect 39117 2363 39175 2369
rect 37967 2329 37979 2332
rect 37921 2323 37979 2329
rect 39117 2329 39129 2363
rect 39163 2360 39175 2363
rect 44376 2360 44404 2391
rect 45094 2388 45100 2440
rect 45152 2428 45158 2440
rect 45373 2431 45431 2437
rect 45373 2428 45385 2431
rect 45152 2400 45385 2428
rect 45152 2388 45158 2400
rect 45373 2397 45385 2400
rect 45419 2397 45431 2431
rect 45373 2391 45431 2397
rect 45922 2388 45928 2440
rect 45980 2428 45986 2440
rect 46201 2431 46259 2437
rect 46201 2428 46213 2431
rect 45980 2400 46213 2428
rect 45980 2388 45986 2400
rect 46201 2397 46213 2400
rect 46247 2397 46259 2431
rect 46201 2391 46259 2397
rect 47029 2431 47087 2437
rect 47029 2397 47041 2431
rect 47075 2428 47087 2431
rect 47486 2428 47492 2440
rect 47075 2400 47492 2428
rect 47075 2397 47087 2400
rect 47029 2391 47087 2397
rect 47486 2388 47492 2400
rect 47544 2388 47550 2440
rect 47581 2431 47639 2437
rect 47581 2397 47593 2431
rect 47627 2397 47639 2431
rect 47762 2428 47768 2440
rect 47723 2400 47768 2428
rect 47581 2391 47639 2397
rect 47596 2360 47624 2391
rect 47762 2388 47768 2400
rect 47820 2388 47826 2440
rect 48314 2388 48320 2440
rect 48372 2428 48378 2440
rect 48593 2431 48651 2437
rect 48593 2428 48605 2431
rect 48372 2400 48605 2428
rect 48372 2388 48378 2400
rect 48593 2397 48605 2400
rect 48639 2397 48651 2431
rect 48593 2391 48651 2397
rect 49605 2431 49663 2437
rect 49605 2397 49617 2431
rect 49651 2428 49663 2431
rect 49878 2428 49884 2440
rect 49651 2400 49884 2428
rect 49651 2397 49663 2400
rect 49605 2391 49663 2397
rect 49878 2388 49884 2400
rect 49936 2388 49942 2440
rect 52196 2437 52224 2468
rect 62666 2456 62672 2468
rect 62724 2456 62730 2508
rect 63052 2505 63080 2536
rect 63405 2533 63417 2567
rect 63451 2564 63463 2567
rect 64046 2564 64052 2576
rect 63451 2536 64052 2564
rect 63451 2533 63463 2536
rect 63405 2527 63463 2533
rect 64046 2524 64052 2536
rect 64104 2524 64110 2576
rect 65794 2564 65800 2576
rect 64156 2536 65800 2564
rect 63037 2499 63095 2505
rect 63037 2465 63049 2499
rect 63083 2465 63095 2499
rect 64156 2496 64184 2536
rect 65794 2524 65800 2536
rect 65852 2524 65858 2576
rect 65981 2567 66039 2573
rect 65981 2533 65993 2567
rect 66027 2564 66039 2567
rect 66254 2564 66260 2576
rect 66027 2536 66260 2564
rect 66027 2533 66039 2536
rect 65981 2527 66039 2533
rect 66254 2524 66260 2536
rect 66312 2524 66318 2576
rect 67269 2567 67327 2573
rect 67269 2564 67281 2567
rect 66456 2536 67281 2564
rect 66456 2505 66484 2536
rect 67269 2533 67281 2536
rect 67315 2533 67327 2567
rect 67269 2527 67327 2533
rect 67542 2524 67548 2576
rect 67600 2564 67606 2576
rect 69477 2567 69535 2573
rect 69477 2564 69489 2567
rect 67600 2536 69489 2564
rect 67600 2524 67606 2536
rect 69477 2533 69489 2536
rect 69523 2533 69535 2567
rect 69937 2567 69995 2573
rect 69937 2564 69949 2567
rect 69477 2527 69535 2533
rect 69676 2536 69949 2564
rect 63037 2459 63095 2465
rect 63236 2468 64184 2496
rect 66441 2499 66499 2505
rect 50985 2431 51043 2437
rect 50985 2397 50997 2431
rect 51031 2428 51043 2431
rect 52181 2431 52239 2437
rect 51031 2400 52132 2428
rect 51031 2397 51043 2400
rect 50985 2391 51043 2397
rect 39163 2332 43208 2360
rect 39163 2329 39175 2332
rect 39117 2323 39175 2329
rect 33686 2292 33692 2304
rect 32631 2264 33692 2292
rect 32631 2261 32643 2264
rect 32585 2255 32643 2261
rect 33686 2252 33692 2264
rect 33744 2252 33750 2304
rect 36354 2252 36360 2304
rect 36412 2292 36418 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 36412 2264 37473 2292
rect 36412 2252 36418 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 38378 2292 38384 2304
rect 38339 2264 38384 2292
rect 37461 2255 37519 2261
rect 38378 2252 38384 2264
rect 38436 2252 38442 2304
rect 39206 2292 39212 2304
rect 39167 2264 39212 2292
rect 39206 2252 39212 2264
rect 39264 2292 39270 2304
rect 40034 2292 40040 2304
rect 39264 2264 40040 2292
rect 39264 2252 39270 2264
rect 40034 2252 40040 2264
rect 40092 2252 40098 2304
rect 40402 2252 40408 2304
rect 40460 2292 40466 2304
rect 40865 2295 40923 2301
rect 40865 2292 40877 2295
rect 40460 2264 40877 2292
rect 40460 2252 40466 2264
rect 40865 2261 40877 2264
rect 40911 2261 40923 2295
rect 43180 2292 43208 2332
rect 44008 2332 44404 2360
rect 45526 2332 47624 2360
rect 47949 2363 48007 2369
rect 44008 2292 44036 2332
rect 43180 2264 44036 2292
rect 40865 2255 40923 2261
rect 44082 2252 44088 2304
rect 44140 2292 44146 2304
rect 44177 2295 44235 2301
rect 44177 2292 44189 2295
rect 44140 2264 44189 2292
rect 44140 2252 44146 2264
rect 44177 2261 44189 2264
rect 44223 2261 44235 2295
rect 44177 2255 44235 2261
rect 45189 2295 45247 2301
rect 45189 2261 45201 2295
rect 45235 2292 45247 2295
rect 45526 2292 45554 2332
rect 47949 2329 47961 2363
rect 47995 2360 48007 2363
rect 50617 2363 50675 2369
rect 50617 2360 50629 2363
rect 47995 2332 50629 2360
rect 47995 2329 48007 2332
rect 47949 2323 48007 2329
rect 50617 2329 50629 2332
rect 50663 2329 50675 2363
rect 52104 2360 52132 2400
rect 52181 2397 52193 2431
rect 52227 2397 52239 2431
rect 52181 2391 52239 2397
rect 52270 2388 52276 2440
rect 52328 2428 52334 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52328 2400 52745 2428
rect 52328 2388 52334 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 52917 2431 52975 2437
rect 52917 2397 52929 2431
rect 52963 2428 52975 2431
rect 53006 2428 53012 2440
rect 52963 2400 53012 2428
rect 52963 2397 52975 2400
rect 52917 2391 52975 2397
rect 53006 2388 53012 2400
rect 53064 2388 53070 2440
rect 53098 2388 53104 2440
rect 53156 2428 53162 2440
rect 53745 2431 53803 2437
rect 53745 2428 53757 2431
rect 53156 2400 53757 2428
rect 53156 2388 53162 2400
rect 53745 2397 53757 2400
rect 53791 2397 53803 2431
rect 54754 2428 54760 2440
rect 54715 2400 54760 2428
rect 53745 2391 53803 2397
rect 54754 2388 54760 2400
rect 54812 2388 54818 2440
rect 55490 2388 55496 2440
rect 55548 2428 55554 2440
rect 55769 2431 55827 2437
rect 55769 2428 55781 2431
rect 55548 2400 55781 2428
rect 55548 2388 55554 2400
rect 55769 2397 55781 2400
rect 55815 2397 55827 2431
rect 55769 2391 55827 2397
rect 56413 2431 56471 2437
rect 56413 2397 56425 2431
rect 56459 2397 56471 2431
rect 56594 2428 56600 2440
rect 56555 2400 56600 2428
rect 56413 2391 56471 2397
rect 53190 2360 53196 2372
rect 52104 2332 53196 2360
rect 50617 2323 50675 2329
rect 53190 2320 53196 2332
rect 53248 2320 53254 2372
rect 46842 2292 46848 2304
rect 45235 2264 45554 2292
rect 46803 2264 46848 2292
rect 45235 2261 45247 2264
rect 45189 2255 45247 2261
rect 46842 2252 46848 2264
rect 46900 2252 46906 2304
rect 51997 2295 52055 2301
rect 51997 2261 52009 2295
rect 52043 2292 52055 2295
rect 53006 2292 53012 2304
rect 52043 2264 53012 2292
rect 52043 2261 52055 2264
rect 51997 2255 52055 2261
rect 53006 2252 53012 2264
rect 53064 2252 53070 2304
rect 54573 2295 54631 2301
rect 54573 2261 54585 2295
rect 54619 2292 54631 2295
rect 56428 2292 56456 2391
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 57882 2388 57888 2440
rect 57940 2428 57946 2440
rect 58161 2431 58219 2437
rect 58161 2428 58173 2431
rect 57940 2400 58173 2428
rect 57940 2388 57946 2400
rect 58161 2397 58173 2400
rect 58207 2397 58219 2431
rect 58161 2391 58219 2397
rect 60366 2388 60372 2440
rect 60424 2428 60430 2440
rect 63236 2437 63264 2468
rect 66441 2465 66453 2499
rect 66487 2465 66499 2499
rect 66806 2496 66812 2508
rect 66767 2468 66812 2496
rect 66441 2459 66499 2465
rect 66806 2456 66812 2468
rect 66864 2456 66870 2508
rect 68830 2496 68836 2508
rect 67606 2468 68692 2496
rect 68791 2468 68836 2496
rect 60645 2431 60703 2437
rect 60645 2428 60657 2431
rect 60424 2400 60657 2428
rect 60424 2388 60430 2400
rect 60645 2397 60657 2400
rect 60691 2397 60703 2431
rect 60645 2391 60703 2397
rect 61657 2431 61715 2437
rect 61657 2397 61669 2431
rect 61703 2397 61715 2431
rect 61657 2391 61715 2397
rect 61749 2431 61807 2437
rect 61749 2397 61761 2431
rect 61795 2428 61807 2431
rect 63221 2431 63279 2437
rect 63221 2428 63233 2431
rect 61795 2400 63233 2428
rect 61795 2397 61807 2400
rect 61749 2391 61807 2397
rect 63221 2397 63233 2400
rect 63267 2397 63279 2431
rect 64049 2431 64107 2437
rect 64049 2428 64061 2431
rect 63221 2391 63279 2397
rect 63604 2400 64061 2428
rect 56781 2363 56839 2369
rect 56781 2329 56793 2363
rect 56827 2360 56839 2363
rect 59541 2363 59599 2369
rect 59541 2360 59553 2363
rect 56827 2332 59553 2360
rect 56827 2329 56839 2332
rect 56781 2323 56839 2329
rect 59541 2329 59553 2332
rect 59587 2329 59599 2363
rect 61672 2360 61700 2391
rect 62114 2360 62120 2372
rect 61672 2332 62120 2360
rect 59541 2323 59599 2329
rect 62114 2320 62120 2332
rect 62172 2320 62178 2372
rect 62758 2320 62764 2372
rect 62816 2360 62822 2372
rect 63604 2360 63632 2400
rect 64049 2397 64061 2400
rect 64095 2397 64107 2431
rect 64049 2391 64107 2397
rect 64322 2388 64328 2440
rect 64380 2428 64386 2440
rect 64693 2431 64751 2437
rect 64693 2428 64705 2431
rect 64380 2400 64705 2428
rect 64380 2388 64386 2400
rect 64693 2397 64705 2400
rect 64739 2397 64751 2431
rect 64693 2391 64751 2397
rect 65613 2431 65671 2437
rect 65613 2397 65625 2431
rect 65659 2397 65671 2431
rect 65794 2428 65800 2440
rect 65755 2400 65800 2428
rect 65613 2391 65671 2397
rect 62816 2332 63632 2360
rect 62816 2320 62822 2332
rect 59814 2292 59820 2304
rect 54619 2264 56456 2292
rect 59775 2264 59820 2292
rect 54619 2261 54631 2264
rect 54573 2255 54631 2261
rect 59814 2252 59820 2264
rect 59872 2252 59878 2304
rect 64509 2295 64567 2301
rect 64509 2261 64521 2295
rect 64555 2292 64567 2295
rect 65628 2292 65656 2391
rect 65794 2388 65800 2400
rect 65852 2428 65858 2440
rect 66625 2431 66683 2437
rect 66625 2428 66637 2431
rect 65852 2400 66637 2428
rect 65852 2388 65858 2400
rect 66625 2397 66637 2400
rect 66671 2397 66683 2431
rect 66625 2391 66683 2397
rect 66640 2360 66668 2391
rect 66714 2388 66720 2440
rect 66772 2428 66778 2440
rect 67453 2431 67511 2437
rect 67453 2428 67465 2431
rect 66772 2400 67465 2428
rect 66772 2388 66778 2400
rect 67453 2397 67465 2400
rect 67499 2397 67511 2431
rect 67453 2391 67511 2397
rect 67606 2360 67634 2468
rect 68664 2440 68692 2468
rect 68830 2456 68836 2468
rect 68888 2456 68894 2508
rect 68557 2431 68615 2437
rect 68557 2397 68569 2431
rect 68603 2397 68615 2431
rect 68557 2391 68615 2397
rect 66640 2332 67634 2360
rect 68572 2360 68600 2391
rect 68646 2388 68652 2440
rect 68704 2428 68710 2440
rect 68704 2400 68749 2428
rect 68704 2388 68710 2400
rect 69676 2360 69704 2536
rect 69937 2533 69949 2536
rect 69983 2533 69995 2567
rect 69937 2527 69995 2533
rect 71593 2567 71651 2573
rect 71593 2533 71605 2567
rect 71639 2564 71651 2567
rect 73706 2564 73712 2576
rect 71639 2536 73384 2564
rect 73667 2536 73712 2564
rect 71639 2533 71651 2536
rect 71593 2527 71651 2533
rect 70026 2456 70032 2508
rect 70084 2496 70090 2508
rect 73356 2505 73384 2536
rect 73706 2524 73712 2536
rect 73764 2524 73770 2576
rect 73816 2536 78996 2564
rect 70949 2499 71007 2505
rect 70949 2496 70961 2499
rect 70084 2468 70961 2496
rect 70084 2456 70090 2468
rect 70949 2465 70961 2468
rect 70995 2465 71007 2499
rect 70949 2459 71007 2465
rect 73341 2499 73399 2505
rect 73341 2465 73353 2499
rect 73387 2465 73399 2499
rect 73816 2496 73844 2536
rect 73341 2459 73399 2465
rect 73448 2468 73844 2496
rect 70118 2428 70124 2440
rect 68572 2332 69704 2360
rect 69860 2400 69980 2428
rect 70079 2400 70124 2428
rect 64555 2264 65656 2292
rect 64555 2261 64567 2264
rect 64509 2255 64567 2261
rect 65702 2252 65708 2304
rect 65760 2292 65766 2304
rect 69860 2292 69888 2400
rect 69952 2360 69980 2400
rect 70118 2388 70124 2400
rect 70176 2388 70182 2440
rect 71498 2388 71504 2440
rect 71556 2428 71562 2440
rect 71777 2431 71835 2437
rect 71777 2428 71789 2431
rect 71556 2400 71789 2428
rect 71556 2388 71562 2400
rect 71777 2397 71789 2400
rect 71823 2397 71835 2431
rect 71777 2391 71835 2397
rect 72326 2388 72332 2440
rect 72384 2428 72390 2440
rect 72605 2431 72663 2437
rect 72605 2428 72617 2431
rect 72384 2400 72617 2428
rect 72384 2388 72390 2400
rect 72605 2397 72617 2400
rect 72651 2397 72663 2431
rect 72605 2391 72663 2397
rect 70762 2360 70768 2372
rect 69952 2332 70768 2360
rect 70762 2320 70768 2332
rect 70820 2360 70826 2372
rect 73448 2360 73476 2468
rect 74534 2456 74540 2508
rect 74592 2496 74598 2508
rect 74592 2468 74637 2496
rect 74592 2456 74598 2468
rect 76374 2456 76380 2508
rect 76432 2496 76438 2508
rect 77021 2499 77079 2505
rect 77021 2496 77033 2499
rect 76432 2468 77033 2496
rect 76432 2456 76438 2468
rect 77021 2465 77033 2468
rect 77067 2465 77079 2499
rect 78968 2496 78996 2536
rect 79042 2524 79048 2576
rect 79100 2564 79106 2576
rect 79962 2564 79968 2576
rect 79100 2536 79968 2564
rect 79100 2524 79106 2536
rect 79962 2524 79968 2536
rect 80020 2564 80026 2576
rect 83093 2567 83151 2573
rect 80020 2536 82952 2564
rect 80020 2524 80026 2536
rect 81986 2496 81992 2508
rect 78968 2468 81992 2496
rect 77021 2459 77079 2465
rect 81986 2456 81992 2468
rect 82044 2456 82050 2508
rect 73525 2431 73583 2437
rect 73525 2397 73537 2431
rect 73571 2428 73583 2431
rect 74721 2431 74779 2437
rect 74721 2428 74733 2431
rect 73571 2400 74733 2428
rect 73571 2397 73583 2400
rect 73525 2391 73583 2397
rect 74721 2397 74733 2400
rect 74767 2397 74779 2431
rect 74721 2391 74779 2397
rect 74905 2431 74963 2437
rect 74905 2397 74917 2431
rect 74951 2428 74963 2431
rect 75917 2431 75975 2437
rect 75917 2428 75929 2431
rect 74951 2400 75929 2428
rect 74951 2397 74963 2400
rect 74905 2391 74963 2397
rect 75917 2397 75929 2400
rect 75963 2397 75975 2431
rect 75917 2391 75975 2397
rect 77205 2431 77263 2437
rect 77205 2397 77217 2431
rect 77251 2397 77263 2431
rect 77205 2391 77263 2397
rect 77389 2431 77447 2437
rect 77389 2397 77401 2431
rect 77435 2428 77447 2431
rect 78493 2431 78551 2437
rect 78493 2428 78505 2431
rect 77435 2400 78505 2428
rect 77435 2397 77447 2400
rect 77389 2391 77447 2397
rect 78493 2397 78505 2400
rect 78539 2397 78551 2431
rect 78493 2391 78551 2397
rect 70820 2332 73476 2360
rect 74736 2360 74764 2391
rect 77220 2360 77248 2391
rect 78674 2388 78680 2440
rect 78732 2428 78738 2440
rect 79413 2431 79471 2437
rect 79413 2428 79425 2431
rect 78732 2400 79425 2428
rect 78732 2388 78738 2400
rect 79413 2397 79425 2400
rect 79459 2397 79471 2431
rect 79413 2391 79471 2397
rect 79502 2388 79508 2440
rect 79560 2428 79566 2440
rect 80057 2431 80115 2437
rect 80057 2428 80069 2431
rect 79560 2400 80069 2428
rect 79560 2388 79566 2400
rect 80057 2397 80069 2400
rect 80103 2397 80115 2431
rect 80057 2391 80115 2397
rect 81342 2388 81348 2440
rect 81400 2428 81406 2440
rect 82096 2437 82124 2536
rect 82924 2437 82952 2536
rect 83093 2533 83105 2567
rect 83139 2564 83151 2567
rect 84856 2564 84884 2604
rect 85390 2592 85396 2604
rect 85448 2592 85454 2644
rect 88150 2632 88156 2644
rect 88111 2604 88156 2632
rect 88150 2592 88156 2604
rect 88208 2592 88214 2644
rect 89438 2632 89444 2644
rect 89399 2604 89444 2632
rect 89438 2592 89444 2604
rect 89496 2592 89502 2644
rect 91741 2635 91799 2641
rect 89686 2604 90588 2632
rect 89686 2564 89714 2604
rect 83139 2536 84792 2564
rect 84856 2536 89714 2564
rect 90560 2564 90588 2604
rect 91741 2601 91753 2635
rect 91787 2632 91799 2635
rect 91830 2632 91836 2644
rect 91787 2604 91836 2632
rect 91787 2601 91799 2604
rect 91741 2595 91799 2601
rect 91830 2592 91836 2604
rect 91888 2592 91894 2644
rect 91922 2592 91928 2644
rect 91980 2632 91986 2644
rect 93213 2635 93271 2641
rect 93213 2632 93225 2635
rect 91980 2604 93225 2632
rect 91980 2592 91986 2604
rect 93213 2601 93225 2604
rect 93259 2601 93271 2635
rect 96890 2632 96896 2644
rect 96851 2604 96896 2632
rect 93213 2595 93271 2601
rect 96890 2592 96896 2604
rect 96948 2592 96954 2644
rect 104986 2632 104992 2644
rect 97000 2604 104992 2632
rect 97000 2564 97028 2604
rect 104986 2592 104992 2604
rect 105044 2592 105050 2644
rect 108298 2632 108304 2644
rect 108259 2604 108304 2632
rect 108298 2592 108304 2604
rect 108356 2592 108362 2644
rect 111061 2635 111119 2641
rect 111061 2601 111073 2635
rect 111107 2632 111119 2635
rect 112254 2632 112260 2644
rect 111107 2604 112260 2632
rect 111107 2601 111119 2604
rect 111061 2595 111119 2601
rect 112254 2592 112260 2604
rect 112312 2592 112318 2644
rect 90560 2536 97028 2564
rect 97721 2567 97779 2573
rect 83139 2533 83151 2536
rect 83093 2527 83151 2533
rect 81437 2431 81495 2437
rect 81437 2428 81449 2431
rect 81400 2400 81449 2428
rect 81400 2388 81406 2400
rect 81437 2397 81449 2400
rect 81483 2397 81495 2431
rect 81437 2391 81495 2397
rect 81897 2431 81955 2437
rect 81897 2397 81909 2431
rect 81943 2397 81955 2431
rect 81897 2391 81955 2397
rect 82081 2431 82139 2437
rect 82081 2397 82093 2431
rect 82127 2397 82139 2431
rect 82725 2431 82783 2437
rect 82725 2428 82737 2431
rect 82081 2391 82139 2397
rect 82188 2400 82737 2428
rect 79042 2360 79048 2372
rect 74736 2332 79048 2360
rect 70820 2320 70826 2332
rect 79042 2320 79048 2332
rect 79100 2320 79106 2372
rect 81912 2360 81940 2391
rect 79244 2332 81940 2360
rect 76098 2292 76104 2304
rect 65760 2264 69888 2292
rect 76059 2264 76104 2292
rect 65760 2252 65766 2264
rect 76098 2252 76104 2264
rect 76156 2252 76162 2304
rect 78677 2295 78735 2301
rect 78677 2261 78689 2295
rect 78723 2292 78735 2295
rect 79134 2292 79140 2304
rect 78723 2264 79140 2292
rect 78723 2261 78735 2264
rect 78677 2255 78735 2261
rect 79134 2252 79140 2264
rect 79192 2252 79198 2304
rect 79244 2301 79272 2332
rect 79229 2295 79287 2301
rect 79229 2261 79241 2295
rect 79275 2261 79287 2295
rect 79229 2255 79287 2261
rect 81253 2295 81311 2301
rect 81253 2261 81265 2295
rect 81299 2292 81311 2295
rect 82188 2292 82216 2400
rect 82725 2397 82737 2400
rect 82771 2397 82783 2431
rect 82725 2391 82783 2397
rect 82909 2431 82967 2437
rect 82909 2397 82921 2431
rect 82955 2397 82967 2431
rect 82909 2391 82967 2397
rect 83550 2388 83556 2440
rect 83608 2428 83614 2440
rect 83829 2431 83887 2437
rect 83829 2428 83841 2431
rect 83608 2400 83841 2428
rect 83608 2388 83614 2400
rect 83829 2397 83841 2400
rect 83875 2397 83887 2431
rect 83829 2391 83887 2397
rect 84286 2388 84292 2440
rect 84344 2428 84350 2440
rect 84565 2431 84623 2437
rect 84565 2428 84577 2431
rect 84344 2400 84577 2428
rect 84344 2388 84350 2400
rect 84565 2397 84577 2400
rect 84611 2397 84623 2431
rect 84764 2428 84792 2536
rect 97721 2533 97733 2567
rect 97767 2564 97779 2567
rect 98086 2564 98092 2576
rect 97767 2536 98092 2564
rect 97767 2533 97779 2536
rect 97721 2527 97779 2533
rect 98086 2524 98092 2536
rect 98144 2524 98150 2576
rect 98181 2567 98239 2573
rect 98181 2533 98193 2567
rect 98227 2533 98239 2567
rect 98181 2527 98239 2533
rect 84838 2456 84844 2508
rect 84896 2496 84902 2508
rect 90450 2496 90456 2508
rect 84896 2468 90456 2496
rect 84896 2456 84902 2468
rect 90450 2456 90456 2468
rect 90508 2456 90514 2508
rect 90652 2468 91600 2496
rect 90652 2440 90680 2468
rect 86681 2431 86739 2437
rect 86681 2428 86693 2431
rect 84764 2400 86693 2428
rect 84565 2391 84623 2397
rect 86681 2397 86693 2400
rect 86727 2397 86739 2431
rect 86681 2391 86739 2397
rect 87877 2431 87935 2437
rect 87877 2397 87889 2431
rect 87923 2397 87935 2431
rect 87877 2391 87935 2397
rect 82265 2363 82323 2369
rect 82265 2329 82277 2363
rect 82311 2360 82323 2363
rect 85301 2363 85359 2369
rect 85301 2360 85313 2363
rect 82311 2332 85313 2360
rect 82311 2329 82323 2332
rect 82265 2323 82323 2329
rect 85301 2329 85313 2332
rect 85347 2329 85359 2363
rect 87892 2360 87920 2391
rect 87966 2388 87972 2440
rect 88024 2428 88030 2440
rect 88024 2400 88069 2428
rect 88024 2388 88030 2400
rect 88150 2388 88156 2440
rect 88208 2428 88214 2440
rect 88981 2431 89039 2437
rect 88981 2428 88993 2431
rect 88208 2400 88993 2428
rect 88208 2388 88214 2400
rect 88981 2397 88993 2400
rect 89027 2397 89039 2431
rect 89622 2428 89628 2440
rect 89583 2400 89628 2428
rect 88981 2391 89039 2397
rect 89622 2388 89628 2400
rect 89680 2388 89686 2440
rect 90542 2428 90548 2440
rect 90503 2400 90548 2428
rect 90542 2388 90548 2400
rect 90600 2388 90606 2440
rect 90634 2388 90640 2440
rect 90692 2428 90698 2440
rect 91572 2437 91600 2468
rect 91646 2456 91652 2508
rect 91704 2496 91710 2508
rect 92569 2499 92627 2505
rect 92569 2496 92581 2499
rect 91704 2468 92581 2496
rect 91704 2456 91710 2468
rect 92569 2465 92581 2468
rect 92615 2465 92627 2499
rect 92569 2459 92627 2465
rect 93946 2456 93952 2508
rect 94004 2496 94010 2508
rect 94777 2499 94835 2505
rect 94777 2496 94789 2499
rect 94004 2468 94789 2496
rect 94004 2456 94010 2468
rect 94777 2465 94789 2468
rect 94823 2465 94835 2499
rect 94777 2459 94835 2465
rect 97353 2499 97411 2505
rect 97353 2465 97365 2499
rect 97399 2496 97411 2499
rect 98196 2496 98224 2527
rect 100294 2524 100300 2576
rect 100352 2564 100358 2576
rect 101861 2567 101919 2573
rect 101861 2564 101873 2567
rect 100352 2536 101873 2564
rect 100352 2524 100358 2536
rect 101861 2533 101873 2536
rect 101907 2533 101919 2567
rect 101861 2527 101919 2533
rect 106001 2567 106059 2573
rect 106001 2533 106013 2567
rect 106047 2564 106059 2567
rect 106047 2536 112300 2564
rect 106047 2533 106059 2536
rect 106001 2527 106059 2533
rect 97399 2468 98224 2496
rect 97399 2465 97411 2468
rect 97353 2459 97411 2465
rect 99006 2456 99012 2508
rect 99064 2496 99070 2508
rect 99101 2499 99159 2505
rect 99101 2496 99113 2499
rect 99064 2468 99113 2496
rect 99064 2456 99070 2468
rect 99101 2465 99113 2468
rect 99147 2465 99159 2499
rect 99101 2459 99159 2465
rect 102318 2456 102324 2508
rect 102376 2496 102382 2508
rect 104621 2499 104679 2505
rect 104621 2496 104633 2499
rect 102376 2468 104633 2496
rect 102376 2456 102382 2468
rect 104621 2465 104633 2468
rect 104667 2465 104679 2499
rect 109954 2496 109960 2508
rect 109915 2468 109960 2496
rect 104621 2459 104679 2465
rect 109954 2456 109960 2468
rect 110012 2496 110018 2508
rect 111613 2499 111671 2505
rect 111613 2496 111625 2499
rect 110012 2468 111625 2496
rect 110012 2456 110018 2468
rect 111613 2465 111625 2468
rect 111659 2465 111671 2499
rect 111613 2459 111671 2465
rect 91373 2431 91431 2437
rect 90692 2400 90737 2428
rect 90692 2388 90698 2400
rect 91373 2397 91385 2431
rect 91419 2397 91431 2431
rect 91373 2391 91431 2397
rect 91557 2431 91615 2437
rect 91557 2397 91569 2431
rect 91603 2397 91615 2431
rect 91557 2391 91615 2397
rect 92293 2431 92351 2437
rect 92293 2397 92305 2431
rect 92339 2397 92351 2431
rect 92293 2391 92351 2397
rect 89438 2360 89444 2372
rect 85301 2323 85359 2329
rect 85408 2332 87828 2360
rect 87892 2332 89444 2360
rect 81299 2264 82216 2292
rect 83645 2295 83703 2301
rect 81299 2261 81311 2264
rect 81253 2255 81311 2261
rect 83645 2261 83657 2295
rect 83691 2292 83703 2295
rect 85408 2292 85436 2332
rect 86770 2292 86776 2304
rect 83691 2264 85436 2292
rect 86731 2264 86776 2292
rect 83691 2261 83703 2264
rect 83645 2255 83703 2261
rect 86770 2252 86776 2264
rect 86828 2252 86834 2304
rect 87800 2292 87828 2332
rect 89438 2320 89444 2332
rect 89496 2320 89502 2372
rect 91388 2360 91416 2391
rect 89686 2332 91416 2360
rect 91572 2360 91600 2391
rect 92308 2360 92336 2391
rect 92382 2388 92388 2440
rect 92440 2428 92446 2440
rect 92440 2400 92485 2428
rect 92440 2388 92446 2400
rect 93394 2388 93400 2440
rect 93452 2428 93458 2440
rect 94133 2431 94191 2437
rect 94133 2428 94145 2431
rect 93452 2400 94145 2428
rect 93452 2388 93458 2400
rect 94133 2397 94145 2400
rect 94179 2397 94191 2431
rect 94133 2391 94191 2397
rect 95510 2388 95516 2440
rect 95568 2428 95574 2440
rect 95789 2431 95847 2437
rect 95789 2428 95801 2431
rect 95568 2400 95801 2428
rect 95568 2388 95574 2400
rect 95789 2397 95801 2400
rect 95835 2397 95847 2431
rect 95789 2391 95847 2397
rect 96525 2431 96583 2437
rect 96525 2397 96537 2431
rect 96571 2397 96583 2431
rect 96706 2428 96712 2440
rect 96667 2400 96712 2428
rect 96525 2391 96583 2397
rect 91572 2332 92244 2360
rect 92308 2332 93992 2360
rect 89686 2292 89714 2332
rect 87800 2264 89714 2292
rect 90821 2295 90879 2301
rect 90821 2261 90833 2295
rect 90867 2292 90879 2295
rect 92014 2292 92020 2304
rect 90867 2264 92020 2292
rect 90867 2261 90879 2264
rect 90821 2255 90879 2261
rect 92014 2252 92020 2264
rect 92072 2252 92078 2304
rect 92216 2292 92244 2332
rect 92382 2292 92388 2304
rect 92216 2264 92388 2292
rect 92382 2252 92388 2264
rect 92440 2252 92446 2304
rect 93964 2301 93992 2332
rect 93949 2295 94007 2301
rect 93949 2261 93961 2295
rect 93995 2261 94007 2295
rect 93949 2255 94007 2261
rect 95605 2295 95663 2301
rect 95605 2261 95617 2295
rect 95651 2292 95663 2295
rect 96540 2292 96568 2391
rect 96706 2388 96712 2400
rect 96764 2428 96770 2440
rect 97537 2431 97595 2437
rect 97537 2428 97549 2431
rect 96764 2400 97549 2428
rect 96764 2388 96770 2400
rect 97537 2397 97549 2400
rect 97583 2397 97595 2431
rect 97537 2391 97595 2397
rect 97902 2388 97908 2440
rect 97960 2428 97966 2440
rect 98365 2431 98423 2437
rect 98365 2428 98377 2431
rect 97960 2400 98377 2428
rect 97960 2388 97966 2400
rect 98365 2397 98377 2400
rect 98411 2397 98423 2431
rect 100938 2428 100944 2440
rect 100899 2400 100944 2428
rect 98365 2391 98423 2397
rect 100938 2388 100944 2400
rect 100996 2388 101002 2440
rect 101677 2431 101735 2437
rect 101677 2428 101689 2431
rect 101232 2400 101689 2428
rect 99368 2363 99426 2369
rect 99368 2329 99380 2363
rect 99414 2360 99426 2363
rect 99414 2332 100800 2360
rect 99414 2329 99426 2332
rect 99368 2323 99426 2329
rect 95651 2264 96568 2292
rect 95651 2261 95663 2264
rect 95605 2255 95663 2261
rect 100386 2252 100392 2304
rect 100444 2292 100450 2304
rect 100772 2301 100800 2332
rect 101232 2304 101260 2400
rect 101677 2397 101689 2400
rect 101723 2428 101735 2431
rect 102229 2431 102287 2437
rect 102229 2428 102241 2431
rect 101723 2400 102241 2428
rect 101723 2397 101735 2400
rect 101677 2391 101735 2397
rect 102229 2397 102241 2400
rect 102275 2397 102287 2431
rect 102778 2428 102784 2440
rect 102739 2400 102784 2428
rect 102229 2391 102287 2397
rect 102778 2388 102784 2400
rect 102836 2428 102842 2440
rect 104894 2437 104900 2440
rect 103333 2431 103391 2437
rect 103333 2428 103345 2431
rect 102836 2400 103345 2428
rect 102836 2388 102842 2400
rect 103333 2397 103345 2400
rect 103379 2428 103391 2431
rect 104888 2428 104900 2437
rect 103379 2400 103514 2428
rect 104855 2400 104900 2428
rect 103379 2397 103391 2400
rect 103333 2391 103391 2397
rect 103486 2360 103514 2400
rect 104888 2391 104900 2400
rect 104894 2388 104900 2391
rect 104952 2388 104958 2440
rect 107562 2428 107568 2440
rect 107523 2400 107568 2428
rect 107562 2388 107568 2400
rect 107620 2388 107626 2440
rect 108485 2431 108543 2437
rect 108485 2397 108497 2431
rect 108531 2428 108543 2431
rect 109770 2428 109776 2440
rect 108531 2400 109448 2428
rect 109731 2400 109776 2428
rect 108531 2397 108543 2400
rect 108485 2391 108543 2397
rect 103793 2363 103851 2369
rect 103793 2360 103805 2363
rect 103486 2332 103805 2360
rect 103793 2329 103805 2332
rect 103839 2360 103851 2363
rect 104437 2363 104495 2369
rect 104437 2360 104449 2363
rect 103839 2332 104449 2360
rect 103839 2329 103851 2332
rect 103793 2323 103851 2329
rect 104437 2329 104449 2332
rect 104483 2329 104495 2363
rect 104437 2323 104495 2329
rect 100481 2295 100539 2301
rect 100481 2292 100493 2295
rect 100444 2264 100493 2292
rect 100444 2252 100450 2264
rect 100481 2261 100493 2264
rect 100527 2261 100539 2295
rect 100481 2255 100539 2261
rect 100757 2295 100815 2301
rect 100757 2261 100769 2295
rect 100803 2261 100815 2295
rect 101214 2292 101220 2304
rect 101175 2264 101220 2292
rect 100757 2255 100815 2261
rect 101214 2252 101220 2264
rect 101272 2252 101278 2304
rect 102686 2252 102692 2304
rect 102744 2292 102750 2304
rect 102965 2295 103023 2301
rect 102965 2292 102977 2295
rect 102744 2264 102977 2292
rect 102744 2252 102750 2264
rect 102965 2261 102977 2264
rect 103011 2261 103023 2295
rect 102965 2255 103023 2261
rect 107470 2252 107476 2304
rect 107528 2292 107534 2304
rect 109420 2301 109448 2400
rect 109770 2388 109776 2400
rect 109828 2388 109834 2440
rect 109862 2388 109868 2440
rect 109920 2428 109926 2440
rect 110785 2431 110843 2437
rect 110785 2428 110797 2431
rect 109920 2400 110797 2428
rect 109920 2388 109926 2400
rect 110785 2397 110797 2400
rect 110831 2397 110843 2431
rect 110785 2391 110843 2397
rect 111429 2431 111487 2437
rect 111429 2397 111441 2431
rect 111475 2428 111487 2431
rect 112070 2428 112076 2440
rect 111475 2400 112076 2428
rect 111475 2397 111487 2400
rect 111429 2391 111487 2397
rect 112070 2388 112076 2400
rect 112128 2388 112134 2440
rect 112165 2431 112223 2437
rect 112165 2397 112177 2431
rect 112211 2397 112223 2431
rect 112165 2391 112223 2397
rect 110690 2320 110696 2372
rect 110748 2360 110754 2372
rect 112180 2360 112208 2391
rect 110748 2332 112208 2360
rect 112272 2360 112300 2536
rect 112346 2524 112352 2576
rect 112404 2564 112410 2576
rect 113361 2567 113419 2573
rect 113361 2564 113373 2567
rect 112404 2536 113373 2564
rect 112404 2524 112410 2536
rect 113361 2533 113373 2536
rect 113407 2533 113419 2567
rect 113361 2527 113419 2533
rect 112806 2388 112812 2440
rect 112864 2428 112870 2440
rect 113177 2431 113235 2437
rect 113177 2428 113189 2431
rect 112864 2400 113189 2428
rect 112864 2388 112870 2400
rect 113177 2397 113189 2400
rect 113223 2397 113235 2431
rect 114554 2428 114560 2440
rect 114515 2400 114560 2428
rect 113177 2391 113235 2397
rect 114554 2388 114560 2400
rect 114612 2388 114618 2440
rect 115474 2388 115480 2440
rect 115532 2428 115538 2440
rect 115569 2431 115627 2437
rect 115569 2428 115581 2431
rect 115532 2400 115581 2428
rect 115532 2388 115538 2400
rect 115569 2397 115581 2400
rect 115615 2397 115627 2431
rect 115842 2428 115848 2440
rect 115803 2400 115848 2428
rect 115569 2391 115627 2397
rect 115842 2388 115848 2400
rect 115900 2388 115906 2440
rect 117130 2428 117136 2440
rect 117091 2400 117136 2428
rect 117130 2388 117136 2400
rect 117188 2388 117194 2440
rect 117222 2388 117228 2440
rect 117280 2428 117286 2440
rect 117869 2431 117927 2437
rect 117869 2428 117881 2431
rect 117280 2400 117881 2428
rect 117280 2388 117286 2400
rect 117869 2397 117881 2400
rect 117915 2397 117927 2431
rect 117869 2391 117927 2397
rect 117406 2360 117412 2372
rect 112272 2332 117412 2360
rect 110748 2320 110754 2332
rect 117406 2320 117412 2332
rect 117464 2320 117470 2372
rect 107749 2295 107807 2301
rect 107749 2292 107761 2295
rect 107528 2264 107761 2292
rect 107528 2252 107534 2264
rect 107749 2261 107761 2264
rect 107795 2261 107807 2295
rect 107749 2255 107807 2261
rect 109405 2295 109463 2301
rect 109405 2261 109417 2295
rect 109451 2261 109463 2295
rect 109405 2255 109463 2261
rect 109865 2295 109923 2301
rect 109865 2261 109877 2295
rect 109911 2292 109923 2295
rect 110601 2295 110659 2301
rect 110601 2292 110613 2295
rect 109911 2264 110613 2292
rect 109911 2261 109923 2264
rect 109865 2255 109923 2261
rect 110601 2261 110613 2264
rect 110647 2261 110659 2295
rect 110601 2255 110659 2261
rect 111521 2295 111579 2301
rect 111521 2261 111533 2295
rect 111567 2292 111579 2295
rect 111981 2295 112039 2301
rect 111981 2292 111993 2295
rect 111567 2264 111993 2292
rect 111567 2261 111579 2264
rect 111521 2255 111579 2261
rect 111981 2261 111993 2264
rect 112027 2261 112039 2295
rect 112806 2292 112812 2304
rect 112767 2264 112812 2292
rect 111981 2255 112039 2261
rect 112806 2252 112812 2264
rect 112864 2252 112870 2304
rect 113910 2252 113916 2304
rect 113968 2292 113974 2304
rect 114741 2295 114799 2301
rect 114741 2292 114753 2295
rect 113968 2264 114753 2292
rect 113968 2252 113974 2264
rect 114741 2261 114753 2264
rect 114787 2261 114799 2295
rect 114741 2255 114799 2261
rect 116302 2252 116308 2304
rect 116360 2292 116366 2304
rect 117317 2295 117375 2301
rect 117317 2292 117329 2295
rect 116360 2264 117329 2292
rect 116360 2252 116366 2264
rect 117317 2261 117329 2264
rect 117363 2261 117375 2295
rect 117317 2255 117375 2261
rect 117866 2252 117872 2304
rect 117924 2292 117930 2304
rect 118053 2295 118111 2301
rect 118053 2292 118065 2295
rect 117924 2264 118065 2292
rect 117924 2252 117930 2264
rect 118053 2261 118065 2264
rect 118099 2261 118111 2295
rect 118053 2255 118111 2261
rect 1104 2202 118864 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 81014 2202
rect 81066 2150 81078 2202
rect 81130 2150 81142 2202
rect 81194 2150 81206 2202
rect 81258 2150 81270 2202
rect 81322 2150 111734 2202
rect 111786 2150 111798 2202
rect 111850 2150 111862 2202
rect 111914 2150 111926 2202
rect 111978 2150 111990 2202
rect 112042 2150 118864 2202
rect 1104 2128 118864 2150
rect 26878 2048 26884 2100
rect 26936 2088 26942 2100
rect 32122 2088 32128 2100
rect 26936 2060 32128 2088
rect 26936 2048 26942 2060
rect 32122 2048 32128 2060
rect 32180 2048 32186 2100
rect 35066 2048 35072 2100
rect 35124 2088 35130 2100
rect 39206 2088 39212 2100
rect 35124 2060 39212 2088
rect 35124 2048 35130 2060
rect 39206 2048 39212 2060
rect 39264 2048 39270 2100
rect 44082 2048 44088 2100
rect 44140 2088 44146 2100
rect 47762 2088 47768 2100
rect 44140 2060 47768 2088
rect 44140 2048 44146 2060
rect 47762 2048 47768 2060
rect 47820 2048 47826 2100
rect 59814 2048 59820 2100
rect 59872 2088 59878 2100
rect 107562 2088 107568 2100
rect 59872 2060 107568 2088
rect 59872 2048 59878 2060
rect 107562 2048 107568 2060
rect 107620 2048 107626 2100
rect 7834 1980 7840 2032
rect 7892 2020 7898 2032
rect 34974 2020 34980 2032
rect 7892 1992 34980 2020
rect 7892 1980 7898 1992
rect 34974 1980 34980 1992
rect 35032 1980 35038 2032
rect 46842 1980 46848 2032
rect 46900 2020 46906 2032
rect 54846 2020 54852 2032
rect 46900 1992 54852 2020
rect 46900 1980 46906 1992
rect 54846 1980 54852 1992
rect 54904 1980 54910 2032
rect 76098 1980 76104 2032
rect 76156 2020 76162 2032
rect 114554 2020 114560 2032
rect 76156 1992 114560 2020
rect 76156 1980 76162 1992
rect 114554 1980 114560 1992
rect 114612 1980 114618 2032
rect 38378 1912 38384 1964
rect 38436 1952 38442 1964
rect 46474 1952 46480 1964
rect 38436 1924 46480 1952
rect 38436 1912 38442 1924
rect 46474 1912 46480 1924
rect 46532 1912 46538 1964
rect 81986 1912 81992 1964
rect 82044 1952 82050 1964
rect 84838 1952 84844 1964
rect 82044 1924 84844 1952
rect 82044 1912 82050 1924
rect 84838 1912 84844 1924
rect 84896 1912 84902 1964
rect 86770 1912 86776 1964
rect 86828 1952 86834 1964
rect 117222 1952 117228 1964
rect 86828 1924 117228 1952
rect 86828 1912 86834 1924
rect 117222 1912 117228 1924
rect 117280 1912 117286 1964
rect 85390 1844 85396 1896
rect 85448 1884 85454 1896
rect 117130 1884 117136 1896
rect 85448 1856 117136 1884
rect 85448 1844 85454 1856
rect 117130 1844 117136 1856
rect 117188 1844 117194 1896
rect 90450 1776 90456 1828
rect 90508 1816 90514 1828
rect 96706 1816 96712 1828
rect 90508 1788 96712 1816
rect 90508 1776 90514 1788
rect 96706 1776 96712 1788
rect 96764 1776 96770 1828
rect 99374 1776 99380 1828
rect 99432 1816 99438 1828
rect 115842 1816 115848 1828
rect 99432 1788 115848 1816
rect 99432 1776 99438 1788
rect 115842 1776 115848 1788
rect 115900 1776 115906 1828
rect 30650 1708 30656 1760
rect 30708 1748 30714 1760
rect 102778 1748 102784 1760
rect 30708 1720 102784 1748
rect 30708 1708 30714 1720
rect 102778 1708 102784 1720
rect 102836 1708 102842 1760
rect 36538 1640 36544 1692
rect 36596 1680 36602 1692
rect 99558 1680 99564 1692
rect 36596 1652 99564 1680
rect 36596 1640 36602 1652
rect 99558 1640 99564 1652
rect 99616 1640 99622 1692
rect 79134 1572 79140 1624
rect 79192 1612 79198 1624
rect 114830 1612 114836 1624
rect 79192 1584 114836 1612
rect 79192 1572 79198 1584
rect 114830 1572 114836 1584
rect 114888 1572 114894 1624
rect 33686 1504 33692 1556
rect 33744 1544 33750 1556
rect 101214 1544 101220 1556
rect 33744 1516 101220 1544
rect 33744 1504 33750 1516
rect 101214 1504 101220 1516
rect 101272 1504 101278 1556
rect 74626 1436 74632 1488
rect 74684 1476 74690 1488
rect 112806 1476 112812 1488
rect 74684 1448 112812 1476
rect 74684 1436 74690 1448
rect 112806 1436 112812 1448
rect 112864 1436 112870 1488
rect 69106 1368 69112 1420
rect 69164 1408 69170 1420
rect 70118 1408 70124 1420
rect 69164 1380 70124 1408
rect 69164 1368 69170 1380
rect 70118 1368 70124 1380
rect 70176 1368 70182 1420
rect 86678 1368 86684 1420
rect 86736 1408 86742 1420
rect 88150 1408 88156 1420
rect 86736 1380 88156 1408
rect 86736 1368 86742 1380
rect 88150 1368 88156 1380
rect 88208 1368 88214 1420
rect 88334 1368 88340 1420
rect 88392 1408 88398 1420
rect 89622 1408 89628 1420
rect 88392 1380 89628 1408
rect 88392 1368 88398 1380
rect 89622 1368 89628 1380
rect 89680 1368 89686 1420
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 96374 37510 96426 37562
rect 96438 37510 96490 37562
rect 96502 37510 96554 37562
rect 96566 37510 96618 37562
rect 96630 37510 96682 37562
rect 1584 37451 1636 37460
rect 1584 37417 1593 37451
rect 1593 37417 1627 37451
rect 1627 37417 1636 37451
rect 1584 37408 1636 37417
rect 2044 37408 2096 37460
rect 14372 37408 14424 37460
rect 22652 37408 22704 37460
rect 26792 37408 26844 37460
rect 30932 37408 30984 37460
rect 35348 37451 35400 37460
rect 35348 37417 35357 37451
rect 35357 37417 35391 37451
rect 35391 37417 35400 37451
rect 35348 37408 35400 37417
rect 86868 37340 86920 37392
rect 50896 37272 50948 37324
rect 76472 37272 76524 37324
rect 92020 37272 92072 37324
rect 10232 37204 10284 37256
rect 39212 37204 39264 37256
rect 47584 37247 47636 37256
rect 47584 37213 47593 37247
rect 47593 37213 47627 37247
rect 47627 37213 47636 37247
rect 47584 37204 47636 37213
rect 51632 37204 51684 37256
rect 54944 37204 54996 37256
rect 59268 37204 59320 37256
rect 64144 37247 64196 37256
rect 64144 37213 64153 37247
rect 64153 37213 64187 37247
rect 64187 37213 64196 37247
rect 64144 37204 64196 37213
rect 68192 37204 68244 37256
rect 74632 37204 74684 37256
rect 84844 37247 84896 37256
rect 84844 37213 84853 37247
rect 84853 37213 84887 37247
rect 84887 37213 84896 37247
rect 84844 37204 84896 37213
rect 93032 37204 93084 37256
rect 109684 37247 109736 37256
rect 109684 37213 109693 37247
rect 109693 37213 109727 37247
rect 109727 37213 109736 37247
rect 109684 37204 109736 37213
rect 40500 37179 40552 37188
rect 40500 37145 40509 37179
rect 40509 37145 40543 37179
rect 40543 37145 40552 37179
rect 40500 37136 40552 37145
rect 47492 37068 47544 37120
rect 55772 37068 55824 37120
rect 59912 37068 59964 37120
rect 64052 37068 64104 37120
rect 64420 37068 64472 37120
rect 84752 37068 84804 37120
rect 109592 37068 109644 37120
rect 117504 37111 117556 37120
rect 117504 37077 117513 37111
rect 117513 37077 117547 37111
rect 117547 37077 117556 37111
rect 117504 37068 117556 37077
rect 117872 37068 117924 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 81014 36966 81066 37018
rect 81078 36966 81130 37018
rect 81142 36966 81194 37018
rect 81206 36966 81258 37018
rect 81270 36966 81322 37018
rect 111734 36966 111786 37018
rect 111798 36966 111850 37018
rect 111862 36966 111914 37018
rect 111926 36966 111978 37018
rect 111990 36966 112042 37018
rect 2780 36864 2832 36916
rect 45560 36864 45612 36916
rect 64144 36864 64196 36916
rect 66352 36864 66404 36916
rect 84844 36864 84896 36916
rect 117228 36864 117280 36916
rect 40500 36796 40552 36848
rect 101772 36796 101824 36848
rect 92112 36728 92164 36780
rect 88708 36524 88760 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 96374 36422 96426 36474
rect 96438 36422 96490 36474
rect 96502 36422 96554 36474
rect 96566 36422 96618 36474
rect 96630 36422 96682 36474
rect 1492 36159 1544 36168
rect 1492 36125 1501 36159
rect 1501 36125 1535 36159
rect 1535 36125 1544 36159
rect 1492 36116 1544 36125
rect 86500 36048 86552 36100
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 81014 35878 81066 35930
rect 81078 35878 81130 35930
rect 81142 35878 81194 35930
rect 81206 35878 81258 35930
rect 81270 35878 81322 35930
rect 111734 35878 111786 35930
rect 111798 35878 111850 35930
rect 111862 35878 111914 35930
rect 111926 35878 111978 35930
rect 111990 35878 112042 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 96374 35334 96426 35386
rect 96438 35334 96490 35386
rect 96502 35334 96554 35386
rect 96566 35334 96618 35386
rect 96630 35334 96682 35386
rect 90272 35028 90324 35080
rect 118056 34935 118108 34944
rect 118056 34901 118065 34935
rect 118065 34901 118099 34935
rect 118099 34901 118108 34935
rect 118056 34892 118108 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 81014 34790 81066 34842
rect 81078 34790 81130 34842
rect 81142 34790 81194 34842
rect 81206 34790 81258 34842
rect 81270 34790 81322 34842
rect 111734 34790 111786 34842
rect 111798 34790 111850 34842
rect 111862 34790 111914 34842
rect 111926 34790 111978 34842
rect 111990 34790 112042 34842
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 1584 34391 1636 34400
rect 1584 34357 1593 34391
rect 1593 34357 1627 34391
rect 1627 34357 1636 34391
rect 1584 34348 1636 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 96374 34246 96426 34298
rect 96438 34246 96490 34298
rect 96502 34246 96554 34298
rect 96566 34246 96618 34298
rect 96630 34246 96682 34298
rect 92480 33804 92532 33856
rect 118056 33847 118108 33856
rect 118056 33813 118065 33847
rect 118065 33813 118099 33847
rect 118099 33813 118108 33847
rect 118056 33804 118108 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 81014 33702 81066 33754
rect 81078 33702 81130 33754
rect 81142 33702 81194 33754
rect 81206 33702 81258 33754
rect 81270 33702 81322 33754
rect 111734 33702 111786 33754
rect 111798 33702 111850 33754
rect 111862 33702 111914 33754
rect 111926 33702 111978 33754
rect 111990 33702 112042 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 96374 33158 96426 33210
rect 96438 33158 96490 33210
rect 96502 33158 96554 33210
rect 96566 33158 96618 33210
rect 96630 33158 96682 33210
rect 1492 32852 1544 32904
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 81014 32614 81066 32666
rect 81078 32614 81130 32666
rect 81142 32614 81194 32666
rect 81206 32614 81258 32666
rect 81270 32614 81322 32666
rect 111734 32614 111786 32666
rect 111798 32614 111850 32666
rect 111862 32614 111914 32666
rect 111926 32614 111978 32666
rect 111990 32614 112042 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 96374 32070 96426 32122
rect 96438 32070 96490 32122
rect 96502 32070 96554 32122
rect 96566 32070 96618 32122
rect 96630 32070 96682 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 81014 31526 81066 31578
rect 81078 31526 81130 31578
rect 81142 31526 81194 31578
rect 81206 31526 81258 31578
rect 81270 31526 81322 31578
rect 111734 31526 111786 31578
rect 111798 31526 111850 31578
rect 111862 31526 111914 31578
rect 111926 31526 111978 31578
rect 111990 31526 112042 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 96374 30982 96426 31034
rect 96438 30982 96490 31034
rect 96502 30982 96554 31034
rect 96566 30982 96618 31034
rect 96630 30982 96682 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 81014 30438 81066 30490
rect 81078 30438 81130 30490
rect 81142 30438 81194 30490
rect 81206 30438 81258 30490
rect 81270 30438 81322 30490
rect 111734 30438 111786 30490
rect 111798 30438 111850 30490
rect 111862 30438 111914 30490
rect 111926 30438 111978 30490
rect 111990 30438 112042 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 96374 29894 96426 29946
rect 96438 29894 96490 29946
rect 96502 29894 96554 29946
rect 96566 29894 96618 29946
rect 96630 29894 96682 29946
rect 2044 29588 2096 29640
rect 117964 29563 118016 29572
rect 117964 29529 117973 29563
rect 117973 29529 118007 29563
rect 118007 29529 118016 29563
rect 117964 29520 118016 29529
rect 1584 29495 1636 29504
rect 1584 29461 1593 29495
rect 1593 29461 1627 29495
rect 1627 29461 1636 29495
rect 1584 29452 1636 29461
rect 112444 29452 112496 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 81014 29350 81066 29402
rect 81078 29350 81130 29402
rect 81142 29350 81194 29402
rect 81206 29350 81258 29402
rect 81270 29350 81322 29402
rect 111734 29350 111786 29402
rect 111798 29350 111850 29402
rect 111862 29350 111914 29402
rect 111926 29350 111978 29402
rect 111990 29350 112042 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 96374 28806 96426 28858
rect 96438 28806 96490 28858
rect 96502 28806 96554 28858
rect 96566 28806 96618 28858
rect 96630 28806 96682 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 81014 28262 81066 28314
rect 81078 28262 81130 28314
rect 81142 28262 81194 28314
rect 81206 28262 81258 28314
rect 81270 28262 81322 28314
rect 111734 28262 111786 28314
rect 111798 28262 111850 28314
rect 111862 28262 111914 28314
rect 111926 28262 111978 28314
rect 111990 28262 112042 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 96374 27718 96426 27770
rect 96438 27718 96490 27770
rect 96502 27718 96554 27770
rect 96566 27718 96618 27770
rect 96630 27718 96682 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 81014 27174 81066 27226
rect 81078 27174 81130 27226
rect 81142 27174 81194 27226
rect 81206 27174 81258 27226
rect 81270 27174 81322 27226
rect 111734 27174 111786 27226
rect 111798 27174 111850 27226
rect 111862 27174 111914 27226
rect 111926 27174 111978 27226
rect 111990 27174 112042 27226
rect 64328 26732 64380 26784
rect 118056 26775 118108 26784
rect 118056 26741 118065 26775
rect 118065 26741 118099 26775
rect 118099 26741 118108 26775
rect 118056 26732 118108 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 96374 26630 96426 26682
rect 96438 26630 96490 26682
rect 96502 26630 96554 26682
rect 96566 26630 96618 26682
rect 96630 26630 96682 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 81014 26086 81066 26138
rect 81078 26086 81130 26138
rect 81142 26086 81194 26138
rect 81206 26086 81258 26138
rect 81270 26086 81322 26138
rect 111734 26086 111786 26138
rect 111798 26086 111850 26138
rect 111862 26086 111914 26138
rect 111926 26086 111978 26138
rect 111990 26086 112042 26138
rect 1400 25984 1452 26036
rect 1768 25984 1820 26036
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 1676 25823 1728 25832
rect 1676 25789 1685 25823
rect 1685 25789 1719 25823
rect 1719 25789 1728 25823
rect 1676 25780 1728 25789
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 96374 25542 96426 25594
rect 96438 25542 96490 25594
rect 96502 25542 96554 25594
rect 96566 25542 96618 25594
rect 96630 25542 96682 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 81014 24998 81066 25050
rect 81078 24998 81130 25050
rect 81142 24998 81194 25050
rect 81206 24998 81258 25050
rect 81270 24998 81322 25050
rect 111734 24998 111786 25050
rect 111798 24998 111850 25050
rect 111862 24998 111914 25050
rect 111926 24998 111978 25050
rect 111990 24998 112042 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 96374 24454 96426 24506
rect 96438 24454 96490 24506
rect 96502 24454 96554 24506
rect 96566 24454 96618 24506
rect 96630 24454 96682 24506
rect 1860 24148 1912 24200
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 81014 23910 81066 23962
rect 81078 23910 81130 23962
rect 81142 23910 81194 23962
rect 81206 23910 81258 23962
rect 81270 23910 81322 23962
rect 111734 23910 111786 23962
rect 111798 23910 111850 23962
rect 111862 23910 111914 23962
rect 111926 23910 111978 23962
rect 111990 23910 112042 23962
rect 54116 23468 54168 23520
rect 118056 23579 118108 23588
rect 118056 23545 118065 23579
rect 118065 23545 118099 23579
rect 118099 23545 118108 23579
rect 118056 23536 118108 23545
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 96374 23366 96426 23418
rect 96438 23366 96490 23418
rect 96502 23366 96554 23418
rect 96566 23366 96618 23418
rect 96630 23366 96682 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 81014 22822 81066 22874
rect 81078 22822 81130 22874
rect 81142 22822 81194 22874
rect 81206 22822 81258 22874
rect 81270 22822 81322 22874
rect 111734 22822 111786 22874
rect 111798 22822 111850 22874
rect 111862 22822 111914 22874
rect 111926 22822 111978 22874
rect 111990 22822 112042 22874
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 68652 22516 68704 22568
rect 52736 22380 52788 22432
rect 118056 22423 118108 22432
rect 118056 22389 118065 22423
rect 118065 22389 118099 22423
rect 118099 22389 118108 22423
rect 118056 22380 118108 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 96374 22278 96426 22330
rect 96438 22278 96490 22330
rect 96502 22278 96554 22330
rect 96566 22278 96618 22330
rect 96630 22278 96682 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 81014 21734 81066 21786
rect 81078 21734 81130 21786
rect 81142 21734 81194 21786
rect 81206 21734 81258 21786
rect 81270 21734 81322 21786
rect 111734 21734 111786 21786
rect 111798 21734 111850 21786
rect 111862 21734 111914 21786
rect 111926 21734 111978 21786
rect 111990 21734 112042 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 96374 21190 96426 21242
rect 96438 21190 96490 21242
rect 96502 21190 96554 21242
rect 96566 21190 96618 21242
rect 96630 21190 96682 21242
rect 117780 20859 117832 20868
rect 117780 20825 117789 20859
rect 117789 20825 117823 20859
rect 117823 20825 117832 20859
rect 117780 20816 117832 20825
rect 77116 20748 77168 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 81014 20646 81066 20698
rect 81078 20646 81130 20698
rect 81142 20646 81194 20698
rect 81206 20646 81258 20698
rect 81270 20646 81322 20698
rect 111734 20646 111786 20698
rect 111798 20646 111850 20698
rect 111862 20646 111914 20698
rect 111926 20646 111978 20698
rect 111990 20646 112042 20698
rect 68652 20587 68704 20596
rect 68652 20553 68661 20587
rect 68661 20553 68695 20587
rect 68695 20553 68704 20587
rect 68652 20544 68704 20553
rect 69296 20544 69348 20596
rect 70400 20544 70452 20596
rect 74632 20587 74684 20596
rect 70676 20476 70728 20528
rect 1676 20340 1728 20392
rect 64972 20272 65024 20324
rect 66168 20408 66220 20460
rect 68836 20408 68888 20460
rect 74632 20553 74641 20587
rect 74641 20553 74675 20587
rect 74675 20553 74684 20587
rect 74632 20544 74684 20553
rect 74908 20408 74960 20460
rect 69296 20340 69348 20392
rect 69388 20383 69440 20392
rect 69388 20349 69397 20383
rect 69397 20349 69431 20383
rect 69431 20349 69440 20383
rect 69388 20340 69440 20349
rect 70400 20340 70452 20392
rect 74724 20383 74776 20392
rect 74724 20349 74733 20383
rect 74733 20349 74767 20383
rect 74767 20349 74776 20383
rect 74724 20340 74776 20349
rect 65432 20247 65484 20256
rect 65432 20213 65441 20247
rect 65441 20213 65475 20247
rect 65475 20213 65484 20247
rect 65432 20204 65484 20213
rect 69020 20204 69072 20256
rect 70032 20204 70084 20256
rect 73620 20204 73672 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 96374 20102 96426 20154
rect 96438 20102 96490 20154
rect 96502 20102 96554 20154
rect 96566 20102 96618 20154
rect 96630 20102 96682 20154
rect 64972 20043 65024 20052
rect 64972 20009 64981 20043
rect 64981 20009 65015 20043
rect 65015 20009 65024 20043
rect 64972 20000 65024 20009
rect 68836 20043 68888 20052
rect 68836 20009 68845 20043
rect 68845 20009 68879 20043
rect 68879 20009 68888 20043
rect 68836 20000 68888 20009
rect 74908 20043 74960 20052
rect 74908 20009 74917 20043
rect 74917 20009 74951 20043
rect 74951 20009 74960 20043
rect 74908 20000 74960 20009
rect 68376 19864 68428 19916
rect 69388 19864 69440 19916
rect 69020 19839 69072 19848
rect 69020 19805 69029 19839
rect 69029 19805 69063 19839
rect 69063 19805 69072 19839
rect 69020 19796 69072 19805
rect 73620 19796 73672 19848
rect 64236 19728 64288 19780
rect 1676 19660 1728 19712
rect 64880 19660 64932 19712
rect 70860 19660 70912 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 81014 19558 81066 19610
rect 81078 19558 81130 19610
rect 81142 19558 81194 19610
rect 81206 19558 81258 19610
rect 81270 19558 81322 19610
rect 111734 19558 111786 19610
rect 111798 19558 111850 19610
rect 111862 19558 111914 19610
rect 111926 19558 111978 19610
rect 111990 19558 112042 19610
rect 64236 19499 64288 19508
rect 64236 19465 64245 19499
rect 64245 19465 64279 19499
rect 64279 19465 64288 19499
rect 64236 19456 64288 19465
rect 64880 19456 64932 19508
rect 1676 19431 1728 19440
rect 1676 19397 1685 19431
rect 1685 19397 1719 19431
rect 1719 19397 1728 19431
rect 1676 19388 1728 19397
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 65432 19320 65484 19372
rect 73896 19456 73948 19508
rect 118056 19499 118108 19508
rect 118056 19465 118065 19499
rect 118065 19465 118099 19499
rect 118099 19465 118108 19499
rect 118056 19456 118108 19465
rect 66168 19295 66220 19304
rect 66168 19261 66177 19295
rect 66177 19261 66211 19295
rect 66211 19261 66220 19295
rect 66168 19252 66220 19261
rect 70032 19320 70084 19372
rect 70860 19363 70912 19372
rect 70860 19329 70869 19363
rect 70869 19329 70903 19363
rect 70903 19329 70912 19363
rect 70860 19320 70912 19329
rect 117872 19363 117924 19372
rect 117872 19329 117881 19363
rect 117881 19329 117915 19363
rect 117915 19329 117924 19363
rect 117872 19320 117924 19329
rect 68376 19295 68428 19304
rect 68376 19261 68385 19295
rect 68385 19261 68419 19295
rect 68419 19261 68428 19295
rect 68376 19252 68428 19261
rect 70676 19159 70728 19168
rect 70676 19125 70685 19159
rect 70685 19125 70719 19159
rect 70719 19125 70728 19159
rect 70676 19116 70728 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 96374 19014 96426 19066
rect 96438 19014 96490 19066
rect 96502 19014 96554 19066
rect 96566 19014 96618 19066
rect 96630 19014 96682 19066
rect 57336 18683 57388 18692
rect 57336 18649 57345 18683
rect 57345 18649 57379 18683
rect 57379 18649 57388 18683
rect 57336 18640 57388 18649
rect 117872 18572 117924 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 81014 18470 81066 18522
rect 81078 18470 81130 18522
rect 81142 18470 81194 18522
rect 81206 18470 81258 18522
rect 81270 18470 81322 18522
rect 111734 18470 111786 18522
rect 111798 18470 111850 18522
rect 111862 18470 111914 18522
rect 111926 18470 111978 18522
rect 111990 18470 112042 18522
rect 117780 18275 117832 18284
rect 117780 18241 117789 18275
rect 117789 18241 117823 18275
rect 117823 18241 117832 18275
rect 117780 18232 117832 18241
rect 117872 18071 117924 18080
rect 117872 18037 117881 18071
rect 117881 18037 117915 18071
rect 117915 18037 117924 18071
rect 117872 18028 117924 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 96374 17926 96426 17978
rect 96438 17926 96490 17978
rect 96502 17926 96554 17978
rect 96566 17926 96618 17978
rect 96630 17926 96682 17978
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 1768 17484 1820 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 81014 17382 81066 17434
rect 81078 17382 81130 17434
rect 81142 17382 81194 17434
rect 81206 17382 81258 17434
rect 81270 17382 81322 17434
rect 111734 17382 111786 17434
rect 111798 17382 111850 17434
rect 111862 17382 111914 17434
rect 111926 17382 111978 17434
rect 111990 17382 112042 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 96374 16838 96426 16890
rect 96438 16838 96490 16890
rect 96502 16838 96554 16890
rect 96566 16838 96618 16890
rect 96630 16838 96682 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 81014 16294 81066 16346
rect 81078 16294 81130 16346
rect 81142 16294 81194 16346
rect 81206 16294 81258 16346
rect 81270 16294 81322 16346
rect 111734 16294 111786 16346
rect 111798 16294 111850 16346
rect 111862 16294 111914 16346
rect 111926 16294 111978 16346
rect 111990 16294 112042 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 96374 15750 96426 15802
rect 96438 15750 96490 15802
rect 96502 15750 96554 15802
rect 96566 15750 96618 15802
rect 96630 15750 96682 15802
rect 117780 15419 117832 15428
rect 117780 15385 117789 15419
rect 117789 15385 117823 15419
rect 117823 15385 117832 15419
rect 117780 15376 117832 15385
rect 70492 15308 70544 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 81014 15206 81066 15258
rect 81078 15206 81130 15258
rect 81142 15206 81194 15258
rect 81206 15206 81258 15258
rect 81270 15206 81322 15258
rect 111734 15206 111786 15258
rect 111798 15206 111850 15258
rect 111862 15206 111914 15258
rect 111926 15206 111978 15258
rect 111990 15206 112042 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 96374 14662 96426 14714
rect 96438 14662 96490 14714
rect 96502 14662 96554 14714
rect 96566 14662 96618 14714
rect 96630 14662 96682 14714
rect 1308 14492 1360 14544
rect 1492 14492 1544 14544
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 81014 14118 81066 14170
rect 81078 14118 81130 14170
rect 81142 14118 81194 14170
rect 81206 14118 81258 14170
rect 81270 14118 81322 14170
rect 111734 14118 111786 14170
rect 111798 14118 111850 14170
rect 111862 14118 111914 14170
rect 111926 14118 111978 14170
rect 111990 14118 112042 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 96374 13574 96426 13626
rect 96438 13574 96490 13626
rect 96502 13574 96554 13626
rect 96566 13574 96618 13626
rect 96630 13574 96682 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 81014 13030 81066 13082
rect 81078 13030 81130 13082
rect 81142 13030 81194 13082
rect 81206 13030 81258 13082
rect 81270 13030 81322 13082
rect 111734 13030 111786 13082
rect 111798 13030 111850 13082
rect 111862 13030 111914 13082
rect 111926 13030 111978 13082
rect 111990 13030 112042 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 96374 12486 96426 12538
rect 96438 12486 96490 12538
rect 96502 12486 96554 12538
rect 96566 12486 96618 12538
rect 96630 12486 96682 12538
rect 117228 12155 117280 12164
rect 117228 12121 117237 12155
rect 117237 12121 117271 12155
rect 117271 12121 117280 12155
rect 117228 12112 117280 12121
rect 39672 12044 39724 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 81014 11942 81066 11994
rect 81078 11942 81130 11994
rect 81142 11942 81194 11994
rect 81206 11942 81258 11994
rect 81270 11942 81322 11994
rect 111734 11942 111786 11994
rect 111798 11942 111850 11994
rect 111862 11942 111914 11994
rect 111926 11942 111978 11994
rect 111990 11942 112042 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 96374 11398 96426 11450
rect 96438 11398 96490 11450
rect 96502 11398 96554 11450
rect 96566 11398 96618 11450
rect 96630 11398 96682 11450
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 7564 11024 7616 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 81014 10854 81066 10906
rect 81078 10854 81130 10906
rect 81142 10854 81194 10906
rect 81206 10854 81258 10906
rect 81270 10854 81322 10906
rect 111734 10854 111786 10906
rect 111798 10854 111850 10906
rect 111862 10854 111914 10906
rect 111926 10854 111978 10906
rect 111990 10854 112042 10906
rect 1860 10684 1912 10736
rect 2044 10684 2096 10736
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 96374 10310 96426 10362
rect 96438 10310 96490 10362
rect 96502 10310 96554 10362
rect 96566 10310 96618 10362
rect 96630 10310 96682 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 81014 9766 81066 9818
rect 81078 9766 81130 9818
rect 81142 9766 81194 9818
rect 81206 9766 81258 9818
rect 81270 9766 81322 9818
rect 111734 9766 111786 9818
rect 111798 9766 111850 9818
rect 111862 9766 111914 9818
rect 111926 9766 111978 9818
rect 111990 9766 112042 9818
rect 22100 9528 22152 9580
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 96374 9222 96426 9274
rect 96438 9222 96490 9274
rect 96502 9222 96554 9274
rect 96566 9222 96618 9274
rect 96630 9222 96682 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 81014 8678 81066 8730
rect 81078 8678 81130 8730
rect 81142 8678 81194 8730
rect 81206 8678 81258 8730
rect 81270 8678 81322 8730
rect 111734 8678 111786 8730
rect 111798 8678 111850 8730
rect 111862 8678 111914 8730
rect 111926 8678 111978 8730
rect 111990 8678 112042 8730
rect 22376 8440 22428 8492
rect 22100 8415 22152 8424
rect 22100 8381 22109 8415
rect 22109 8381 22143 8415
rect 22143 8381 22152 8415
rect 22100 8372 22152 8381
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 96374 8134 96426 8186
rect 96438 8134 96490 8186
rect 96502 8134 96554 8186
rect 96566 8134 96618 8186
rect 96630 8134 96682 8186
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 10324 7692 10376 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 81014 7590 81066 7642
rect 81078 7590 81130 7642
rect 81142 7590 81194 7642
rect 81206 7590 81258 7642
rect 81270 7590 81322 7642
rect 111734 7590 111786 7642
rect 111798 7590 111850 7642
rect 111862 7590 111914 7642
rect 111926 7590 111978 7642
rect 111990 7590 112042 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 117964 6715 118016 6724
rect 117964 6681 117973 6715
rect 117973 6681 118007 6715
rect 118007 6681 118016 6715
rect 117964 6672 118016 6681
rect 114468 6604 114520 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 81014 6502 81066 6554
rect 81078 6502 81130 6554
rect 81142 6502 81194 6554
rect 81206 6502 81258 6554
rect 81270 6502 81322 6554
rect 111734 6502 111786 6554
rect 111798 6502 111850 6554
rect 111862 6502 111914 6554
rect 111926 6502 111978 6554
rect 111990 6502 112042 6554
rect 77116 6443 77168 6452
rect 77116 6409 77125 6443
rect 77125 6409 77159 6443
rect 77159 6409 77168 6443
rect 77116 6400 77168 6409
rect 76932 6264 76984 6316
rect 77208 6239 77260 6248
rect 77208 6205 77217 6239
rect 77217 6205 77251 6239
rect 77251 6205 77260 6239
rect 77208 6196 77260 6205
rect 76012 6060 76064 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 75920 5695 75972 5704
rect 75920 5661 75929 5695
rect 75929 5661 75963 5695
rect 75963 5661 75972 5695
rect 75920 5652 75972 5661
rect 76012 5652 76064 5704
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 17132 5516 17184 5568
rect 76932 5516 76984 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 81014 5414 81066 5466
rect 81078 5414 81130 5466
rect 81142 5414 81194 5466
rect 81206 5414 81258 5466
rect 81270 5414 81322 5466
rect 111734 5414 111786 5466
rect 111798 5414 111850 5466
rect 111862 5414 111914 5466
rect 111926 5414 111978 5466
rect 111990 5414 112042 5466
rect 10048 5312 10100 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 17224 5312 17276 5364
rect 20812 5312 20864 5364
rect 39672 5355 39724 5364
rect 7564 5244 7616 5296
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 18420 5176 18472 5228
rect 22192 5219 22244 5228
rect 1952 5040 2004 5092
rect 22192 5185 22201 5219
rect 22201 5185 22235 5219
rect 22235 5185 22244 5219
rect 22192 5176 22244 5185
rect 28632 5219 28684 5228
rect 28632 5185 28641 5219
rect 28641 5185 28675 5219
rect 28675 5185 28684 5219
rect 28632 5176 28684 5185
rect 39672 5321 39681 5355
rect 39681 5321 39715 5355
rect 39715 5321 39724 5355
rect 39672 5312 39724 5321
rect 39856 5312 39908 5364
rect 49884 5312 49936 5364
rect 49976 5355 50028 5364
rect 49976 5321 49985 5355
rect 49985 5321 50019 5355
rect 50019 5321 50028 5355
rect 49976 5312 50028 5321
rect 50068 5312 50120 5364
rect 50896 5355 50948 5364
rect 50896 5321 50905 5355
rect 50905 5321 50939 5355
rect 50939 5321 50948 5355
rect 50896 5312 50948 5321
rect 64420 5355 64472 5364
rect 39580 5219 39632 5228
rect 39580 5185 39589 5219
rect 39589 5185 39623 5219
rect 39623 5185 39632 5219
rect 39580 5176 39632 5185
rect 1768 4972 1820 5024
rect 20812 4972 20864 5024
rect 21364 4972 21416 5024
rect 49332 5176 49384 5228
rect 39856 5151 39908 5160
rect 39856 5117 39865 5151
rect 39865 5117 39899 5151
rect 39899 5117 39908 5151
rect 39856 5108 39908 5117
rect 48596 5151 48648 5160
rect 48596 5117 48605 5151
rect 48605 5117 48639 5151
rect 48639 5117 48648 5151
rect 48596 5108 48648 5117
rect 49884 5108 49936 5160
rect 50988 5151 51040 5160
rect 50988 5117 50997 5151
rect 50997 5117 51031 5151
rect 51031 5117 51040 5151
rect 50988 5108 51040 5117
rect 53564 5219 53616 5228
rect 53564 5185 53573 5219
rect 53573 5185 53607 5219
rect 53607 5185 53616 5219
rect 53564 5176 53616 5185
rect 64420 5321 64429 5355
rect 64429 5321 64463 5355
rect 64463 5321 64472 5355
rect 64420 5312 64472 5321
rect 70492 5355 70544 5364
rect 64052 5176 64104 5228
rect 70492 5321 70501 5355
rect 70501 5321 70535 5355
rect 70535 5321 70544 5355
rect 70492 5312 70544 5321
rect 70124 5176 70176 5228
rect 92020 5355 92072 5364
rect 92020 5321 92029 5355
rect 92029 5321 92063 5355
rect 92063 5321 92072 5355
rect 92020 5312 92072 5321
rect 97632 5312 97684 5364
rect 103796 5312 103848 5364
rect 74448 5244 74500 5296
rect 91928 5219 91980 5228
rect 91928 5185 91937 5219
rect 91937 5185 91971 5219
rect 91971 5185 91980 5219
rect 91928 5176 91980 5185
rect 29736 4972 29788 5024
rect 38660 4972 38712 5024
rect 48596 4972 48648 5024
rect 61660 5040 61712 5092
rect 77208 5108 77260 5160
rect 77300 5040 77352 5092
rect 94044 5108 94096 5160
rect 96804 5176 96856 5228
rect 96988 5219 97040 5228
rect 96988 5185 97022 5219
rect 97022 5185 97040 5219
rect 100760 5219 100812 5228
rect 96988 5176 97040 5185
rect 100760 5185 100769 5219
rect 100769 5185 100803 5219
rect 100803 5185 100812 5219
rect 100760 5176 100812 5185
rect 100300 5151 100352 5160
rect 100300 5117 100309 5151
rect 100309 5117 100343 5151
rect 100343 5117 100352 5151
rect 100300 5108 100352 5117
rect 117780 5244 117832 5296
rect 104532 5176 104584 5228
rect 102324 5151 102376 5160
rect 102324 5117 102333 5151
rect 102333 5117 102367 5151
rect 102367 5117 102376 5151
rect 102324 5108 102376 5117
rect 106464 5151 106516 5160
rect 106464 5117 106473 5151
rect 106473 5117 106507 5151
rect 106507 5117 106516 5151
rect 106464 5108 106516 5117
rect 96620 5040 96672 5092
rect 50068 4972 50120 5024
rect 63040 5015 63092 5024
rect 63040 4981 63049 5015
rect 63049 4981 63083 5015
rect 63083 4981 63092 5015
rect 63040 4972 63092 4981
rect 68560 5015 68612 5024
rect 68560 4981 68569 5015
rect 68569 4981 68603 5015
rect 68603 4981 68612 5015
rect 68560 4972 68612 4981
rect 73436 5015 73488 5024
rect 73436 4981 73445 5015
rect 73445 4981 73479 5015
rect 73479 4981 73488 5015
rect 73436 4972 73488 4981
rect 91100 4972 91152 5024
rect 93952 4972 94004 5024
rect 100208 4972 100260 5024
rect 100944 4972 100996 5024
rect 103796 4972 103848 5024
rect 114468 5040 114520 5092
rect 107844 5015 107896 5024
rect 107844 4981 107853 5015
rect 107853 4981 107887 5015
rect 107887 4981 107896 5015
rect 118056 5015 118108 5024
rect 107844 4972 107896 4981
rect 118056 4981 118065 5015
rect 118065 4981 118099 5015
rect 118099 4981 118108 5015
rect 118056 4972 118108 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 22192 4768 22244 4820
rect 22744 4768 22796 4820
rect 38568 4768 38620 4820
rect 48596 4768 48648 4820
rect 49332 4811 49384 4820
rect 49332 4777 49341 4811
rect 49341 4777 49375 4811
rect 49375 4777 49384 4811
rect 49332 4768 49384 4777
rect 63132 4768 63184 4820
rect 64052 4768 64104 4820
rect 69204 4811 69256 4820
rect 69204 4777 69213 4811
rect 69213 4777 69247 4811
rect 69247 4777 69256 4811
rect 69204 4768 69256 4777
rect 70124 4768 70176 4820
rect 76932 4811 76984 4820
rect 76932 4777 76941 4811
rect 76941 4777 76975 4811
rect 76975 4777 76984 4811
rect 76932 4768 76984 4777
rect 91928 4768 91980 4820
rect 96988 4768 97040 4820
rect 100760 4768 100812 4820
rect 104532 4811 104584 4820
rect 104532 4777 104541 4811
rect 104541 4777 104575 4811
rect 104575 4777 104584 4811
rect 104532 4768 104584 4777
rect 75920 4700 75972 4752
rect 86224 4700 86276 4752
rect 2412 4564 2464 4616
rect 9864 4539 9916 4548
rect 9864 4505 9898 4539
rect 9898 4505 9916 4539
rect 9864 4496 9916 4505
rect 17132 4564 17184 4616
rect 21364 4564 21416 4616
rect 49976 4632 50028 4684
rect 50988 4632 51040 4684
rect 61660 4675 61712 4684
rect 61660 4641 61669 4675
rect 61669 4641 61703 4675
rect 61703 4641 61712 4675
rect 61660 4632 61712 4641
rect 73988 4632 74040 4684
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 50068 4564 50120 4616
rect 50620 4564 50672 4616
rect 53564 4564 53616 4616
rect 63040 4564 63092 4616
rect 68560 4564 68612 4616
rect 10232 4428 10284 4480
rect 28172 4428 28224 4480
rect 28632 4428 28684 4480
rect 69388 4496 69440 4548
rect 73436 4564 73488 4616
rect 93952 4607 94004 4616
rect 75920 4496 75972 4548
rect 76748 4496 76800 4548
rect 50160 4428 50212 4480
rect 73896 4428 73948 4480
rect 74448 4428 74500 4480
rect 90364 4496 90416 4548
rect 93952 4573 93961 4607
rect 93961 4573 93995 4607
rect 93995 4573 94004 4607
rect 93952 4564 94004 4573
rect 94688 4564 94740 4616
rect 100300 4700 100352 4752
rect 105084 4700 105136 4752
rect 109960 4700 110012 4752
rect 97632 4675 97684 4684
rect 97632 4641 97641 4675
rect 97641 4641 97675 4675
rect 97675 4641 97684 4675
rect 97632 4632 97684 4641
rect 107844 4632 107896 4684
rect 112444 4675 112496 4684
rect 112444 4641 112453 4675
rect 112453 4641 112487 4675
rect 112487 4641 112496 4675
rect 112444 4632 112496 4641
rect 100208 4607 100260 4616
rect 94044 4496 94096 4548
rect 94320 4539 94372 4548
rect 94320 4505 94329 4539
rect 94329 4505 94363 4539
rect 94363 4505 94372 4539
rect 94320 4496 94372 4505
rect 94596 4496 94648 4548
rect 100208 4573 100217 4607
rect 100217 4573 100251 4607
rect 100251 4573 100260 4607
rect 100208 4564 100260 4573
rect 100944 4564 100996 4616
rect 104716 4607 104768 4616
rect 104716 4573 104725 4607
rect 104725 4573 104759 4607
rect 104759 4573 104768 4607
rect 104716 4564 104768 4573
rect 107384 4607 107436 4616
rect 107384 4573 107393 4607
rect 107393 4573 107427 4607
rect 107427 4573 107436 4607
rect 107384 4564 107436 4573
rect 100484 4496 100536 4548
rect 78588 4428 78640 4480
rect 96804 4428 96856 4480
rect 99012 4428 99064 4480
rect 102324 4428 102376 4480
rect 106464 4428 106516 4480
rect 107016 4428 107068 4480
rect 107200 4471 107252 4480
rect 107200 4437 107209 4471
rect 107209 4437 107243 4471
rect 107243 4437 107252 4471
rect 107200 4428 107252 4437
rect 111156 4471 111208 4480
rect 111156 4437 111165 4471
rect 111165 4437 111199 4471
rect 111199 4437 111208 4471
rect 111156 4428 111208 4437
rect 112352 4471 112404 4480
rect 112352 4437 112361 4471
rect 112361 4437 112395 4471
rect 112395 4437 112404 4471
rect 112352 4428 112404 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 81014 4326 81066 4378
rect 81078 4326 81130 4378
rect 81142 4326 81194 4378
rect 81206 4326 81258 4378
rect 81270 4326 81322 4378
rect 111734 4326 111786 4378
rect 111798 4326 111850 4378
rect 111862 4326 111914 4378
rect 111926 4326 111978 4378
rect 111990 4326 112042 4378
rect 38752 4224 38804 4276
rect 39580 4224 39632 4276
rect 53564 4224 53616 4276
rect 77300 4224 77352 4276
rect 86316 4224 86368 4276
rect 90364 4267 90416 4276
rect 90364 4233 90373 4267
rect 90373 4233 90407 4267
rect 90407 4233 90416 4267
rect 90364 4224 90416 4233
rect 1400 4088 1452 4140
rect 2596 4088 2648 4140
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 18420 4088 18472 4140
rect 38660 4088 38712 4140
rect 73896 4131 73948 4140
rect 73896 4097 73905 4131
rect 73905 4097 73939 4131
rect 73939 4097 73948 4131
rect 73896 4088 73948 4097
rect 73988 4131 74040 4140
rect 73988 4097 73997 4131
rect 73997 4097 74031 4131
rect 74031 4097 74040 4131
rect 77300 4131 77352 4140
rect 73988 4088 74040 4097
rect 77300 4097 77309 4131
rect 77309 4097 77343 4131
rect 77343 4097 77352 4131
rect 77300 4088 77352 4097
rect 86316 4088 86368 4140
rect 87604 4088 87656 4140
rect 91100 4088 91152 4140
rect 94320 4156 94372 4208
rect 96712 4156 96764 4208
rect 97172 4156 97224 4208
rect 100944 4224 100996 4276
rect 101128 4224 101180 4276
rect 104716 4224 104768 4276
rect 112352 4224 112404 4276
rect 101312 4199 101364 4208
rect 97264 4131 97316 4140
rect 22744 4063 22796 4072
rect 22744 4029 22753 4063
rect 22753 4029 22787 4063
rect 22787 4029 22796 4063
rect 22744 4020 22796 4029
rect 28172 4063 28224 4072
rect 28172 4029 28181 4063
rect 28181 4029 28215 4063
rect 28215 4029 28224 4063
rect 28172 4020 28224 4029
rect 38568 4063 38620 4072
rect 38568 4029 38577 4063
rect 38577 4029 38611 4063
rect 38611 4029 38620 4063
rect 38568 4020 38620 4029
rect 45468 4020 45520 4072
rect 50620 4020 50672 4072
rect 59452 4020 59504 4072
rect 63132 4020 63184 4072
rect 69204 4020 69256 4072
rect 74724 4020 74776 4072
rect 86500 4063 86552 4072
rect 35348 3952 35400 4004
rect 10140 3884 10192 3936
rect 19984 3884 20036 3936
rect 23756 3884 23808 3936
rect 28540 3927 28592 3936
rect 28540 3893 28549 3927
rect 28549 3893 28583 3927
rect 28583 3893 28592 3927
rect 28540 3884 28592 3893
rect 31668 3884 31720 3936
rect 68376 3952 68428 4004
rect 86500 4029 86509 4063
rect 86509 4029 86543 4063
rect 86543 4029 86552 4063
rect 86500 4020 86552 4029
rect 87236 3952 87288 4004
rect 42892 3884 42944 3936
rect 47676 3884 47728 3936
rect 52460 3884 52512 3936
rect 57980 3884 58032 3936
rect 62212 3884 62264 3936
rect 68192 3884 68244 3936
rect 73620 3884 73672 3936
rect 86316 3884 86368 3936
rect 86500 3884 86552 3936
rect 90732 4020 90784 4072
rect 97264 4097 97273 4131
rect 97273 4097 97307 4131
rect 97307 4097 97316 4131
rect 97264 4088 97316 4097
rect 93860 4020 93912 4072
rect 94596 4020 94648 4072
rect 94688 4020 94740 4072
rect 100484 4131 100536 4140
rect 100484 4097 100493 4131
rect 100493 4097 100527 4131
rect 100527 4097 100536 4131
rect 100484 4088 100536 4097
rect 100392 4020 100444 4072
rect 101312 4165 101321 4199
rect 101321 4165 101355 4199
rect 101355 4165 101364 4199
rect 101312 4156 101364 4165
rect 101128 4131 101180 4140
rect 101128 4097 101137 4131
rect 101137 4097 101171 4131
rect 101171 4097 101180 4131
rect 101496 4131 101548 4140
rect 101128 4088 101180 4097
rect 101496 4097 101505 4131
rect 101505 4097 101539 4131
rect 101539 4097 101548 4131
rect 101496 4088 101548 4097
rect 101772 4131 101824 4140
rect 101772 4097 101781 4131
rect 101781 4097 101815 4131
rect 101815 4097 101824 4131
rect 101772 4088 101824 4097
rect 105084 4131 105136 4140
rect 89076 3884 89128 3936
rect 90548 3884 90600 3936
rect 91652 3952 91704 4004
rect 101680 4020 101732 4072
rect 105084 4097 105093 4131
rect 105093 4097 105127 4131
rect 105127 4097 105136 4131
rect 105084 4088 105136 4097
rect 107200 4156 107252 4208
rect 111156 4156 111208 4208
rect 117964 4199 118016 4208
rect 117964 4165 117973 4199
rect 117973 4165 118007 4199
rect 118007 4165 118016 4199
rect 117964 4156 118016 4165
rect 107108 4063 107160 4072
rect 107108 4029 107117 4063
rect 107117 4029 107151 4063
rect 107151 4029 107160 4063
rect 107108 4020 107160 4029
rect 98000 3884 98052 3936
rect 103612 3884 103664 3936
rect 104900 3927 104952 3936
rect 104900 3893 104909 3927
rect 104909 3893 104943 3927
rect 104943 3893 104952 3927
rect 104900 3884 104952 3893
rect 105176 3884 105228 3936
rect 109684 3952 109736 4004
rect 108488 3927 108540 3936
rect 108488 3893 108497 3927
rect 108497 3893 108531 3927
rect 108531 3893 108540 3927
rect 108488 3884 108540 3893
rect 110972 3884 111024 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 2872 3680 2924 3732
rect 59268 3723 59320 3732
rect 35348 3612 35400 3664
rect 38384 3612 38436 3664
rect 45468 3612 45520 3664
rect 45652 3655 45704 3664
rect 45652 3621 45661 3655
rect 45661 3621 45695 3655
rect 45695 3621 45704 3655
rect 45652 3612 45704 3621
rect 47584 3612 47636 3664
rect 47676 3612 47728 3664
rect 52460 3612 52512 3664
rect 59268 3689 59277 3723
rect 59277 3689 59311 3723
rect 59311 3689 59320 3723
rect 59268 3680 59320 3689
rect 79140 3680 79192 3732
rect 1676 3544 1728 3596
rect 52736 3587 52788 3596
rect 52736 3553 52745 3587
rect 52745 3553 52779 3587
rect 52779 3553 52788 3587
rect 52736 3544 52788 3553
rect 54116 3587 54168 3596
rect 54116 3553 54125 3587
rect 54125 3553 54159 3587
rect 54159 3553 54168 3587
rect 54116 3544 54168 3553
rect 59452 3612 59504 3664
rect 73988 3612 74040 3664
rect 87236 3680 87288 3732
rect 91560 3680 91612 3732
rect 91744 3723 91796 3732
rect 91744 3689 91753 3723
rect 91753 3689 91787 3723
rect 91787 3689 91796 3723
rect 91744 3680 91796 3689
rect 92480 3723 92532 3732
rect 92480 3689 92489 3723
rect 92489 3689 92523 3723
rect 92523 3689 92532 3723
rect 92480 3680 92532 3689
rect 98000 3723 98052 3732
rect 98000 3689 98009 3723
rect 98009 3689 98043 3723
rect 98043 3689 98052 3723
rect 98000 3680 98052 3689
rect 100300 3680 100352 3732
rect 107384 3680 107436 3732
rect 109776 3680 109828 3732
rect 94688 3612 94740 3664
rect 117504 3680 117556 3732
rect 64328 3587 64380 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 2596 3476 2648 3528
rect 10140 3519 10192 3528
rect 1952 3408 2004 3460
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 19984 3519 20036 3528
rect 19984 3485 19993 3519
rect 19993 3485 20027 3519
rect 20027 3485 20036 3519
rect 19984 3476 20036 3485
rect 23756 3519 23808 3528
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 38476 3519 38528 3528
rect 37832 3451 37884 3460
rect 388 3340 440 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 10048 3340 10100 3392
rect 19432 3340 19484 3392
rect 24400 3340 24452 3392
rect 28448 3340 28500 3392
rect 37832 3417 37841 3451
rect 37841 3417 37875 3451
rect 37875 3417 37884 3451
rect 37832 3408 37884 3417
rect 38476 3485 38485 3519
rect 38485 3485 38519 3519
rect 38519 3485 38528 3519
rect 38476 3476 38528 3485
rect 38568 3519 38620 3528
rect 38568 3485 38597 3519
rect 38597 3485 38620 3519
rect 38568 3476 38620 3485
rect 42892 3476 42944 3528
rect 45468 3519 45520 3528
rect 45468 3485 45477 3519
rect 45477 3485 45511 3519
rect 45511 3485 45520 3519
rect 45468 3476 45520 3485
rect 40684 3408 40736 3460
rect 46112 3408 46164 3460
rect 40224 3340 40276 3392
rect 46480 3476 46532 3528
rect 47584 3519 47636 3528
rect 47584 3485 47593 3519
rect 47593 3485 47627 3519
rect 47627 3485 47636 3519
rect 47584 3476 47636 3485
rect 50160 3519 50212 3528
rect 50160 3485 50169 3519
rect 50169 3485 50203 3519
rect 50203 3485 50212 3519
rect 50160 3476 50212 3485
rect 52460 3519 52512 3528
rect 52460 3485 52469 3519
rect 52469 3485 52503 3519
rect 52503 3485 52512 3519
rect 52460 3476 52512 3485
rect 52828 3476 52880 3528
rect 46388 3340 46440 3392
rect 53288 3408 53340 3460
rect 56968 3476 57020 3528
rect 64328 3553 64337 3587
rect 64337 3553 64371 3587
rect 64371 3553 64380 3587
rect 64328 3544 64380 3553
rect 78588 3544 78640 3596
rect 86224 3587 86276 3596
rect 86224 3553 86233 3587
rect 86233 3553 86267 3587
rect 86267 3553 86276 3587
rect 86224 3544 86276 3553
rect 87604 3544 87656 3596
rect 91744 3544 91796 3596
rect 91928 3587 91980 3596
rect 91928 3553 91937 3587
rect 91937 3553 91971 3587
rect 91971 3553 91980 3587
rect 91928 3544 91980 3553
rect 93952 3587 94004 3596
rect 93952 3553 93961 3587
rect 93961 3553 93995 3587
rect 93995 3553 94004 3587
rect 93952 3544 94004 3553
rect 97172 3587 97224 3596
rect 97172 3553 97181 3587
rect 97181 3553 97215 3587
rect 97215 3553 97224 3587
rect 97172 3544 97224 3553
rect 62212 3519 62264 3528
rect 62212 3485 62221 3519
rect 62221 3485 62255 3519
rect 62255 3485 62264 3519
rect 62212 3476 62264 3485
rect 64052 3519 64104 3528
rect 64052 3485 64061 3519
rect 64061 3485 64095 3519
rect 64095 3485 64104 3519
rect 64052 3476 64104 3485
rect 66812 3476 66864 3528
rect 68836 3476 68888 3528
rect 73896 3476 73948 3528
rect 83556 3519 83608 3528
rect 83556 3485 83565 3519
rect 83565 3485 83599 3519
rect 83599 3485 83608 3519
rect 83556 3476 83608 3485
rect 86316 3476 86368 3528
rect 61752 3340 61804 3392
rect 62396 3340 62448 3392
rect 74540 3340 74592 3392
rect 83648 3340 83700 3392
rect 88708 3519 88760 3528
rect 88708 3485 88717 3519
rect 88717 3485 88751 3519
rect 88751 3485 88760 3519
rect 88708 3476 88760 3485
rect 87696 3408 87748 3460
rect 91652 3476 91704 3528
rect 95056 3476 95108 3528
rect 91744 3451 91796 3460
rect 91744 3417 91753 3451
rect 91753 3417 91787 3451
rect 91787 3417 91796 3451
rect 91744 3408 91796 3417
rect 91836 3408 91888 3460
rect 89628 3340 89680 3392
rect 91192 3340 91244 3392
rect 94964 3383 95016 3392
rect 94964 3349 94973 3383
rect 94973 3349 95007 3383
rect 95007 3349 95016 3383
rect 94964 3340 95016 3349
rect 99288 3476 99340 3528
rect 101312 3544 101364 3596
rect 101680 3587 101732 3596
rect 101680 3553 101689 3587
rect 101689 3553 101723 3587
rect 101723 3553 101732 3587
rect 101680 3544 101732 3553
rect 101772 3544 101824 3596
rect 103612 3544 103664 3596
rect 100392 3476 100444 3528
rect 101496 3476 101548 3528
rect 97264 3408 97316 3460
rect 96988 3383 97040 3392
rect 96988 3349 96997 3383
rect 96997 3349 97031 3383
rect 97031 3349 97040 3383
rect 96988 3340 97040 3349
rect 98184 3408 98236 3460
rect 108488 3544 108540 3596
rect 108396 3476 108448 3528
rect 111984 3451 112036 3460
rect 100760 3340 100812 3392
rect 111984 3417 111993 3451
rect 111993 3417 112027 3451
rect 112027 3417 112036 3451
rect 111984 3408 112036 3417
rect 112352 3408 112404 3460
rect 115572 3476 115624 3528
rect 117412 3476 117464 3528
rect 112628 3383 112680 3392
rect 112628 3349 112637 3383
rect 112637 3349 112671 3383
rect 112671 3349 112680 3383
rect 112628 3340 112680 3349
rect 118148 3340 118200 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 81014 3238 81066 3290
rect 81078 3238 81130 3290
rect 81142 3238 81194 3290
rect 81206 3238 81258 3290
rect 81270 3238 81322 3290
rect 111734 3238 111786 3290
rect 111798 3238 111850 3290
rect 111862 3238 111914 3290
rect 111926 3238 111978 3290
rect 111990 3238 112042 3290
rect 1400 3136 1452 3188
rect 1492 3068 1544 3120
rect 46204 3136 46256 3188
rect 51908 3136 51960 3188
rect 53288 3179 53340 3188
rect 2228 3000 2280 3052
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 5264 3000 5316 3052
rect 21916 3000 21968 3052
rect 28448 3043 28500 3052
rect 28448 3009 28457 3043
rect 28457 3009 28491 3043
rect 28491 3009 28500 3043
rect 28448 3000 28500 3009
rect 30840 3000 30892 3052
rect 33048 3000 33100 3052
rect 34704 3000 34756 3052
rect 8300 2932 8352 2984
rect 32128 2975 32180 2984
rect 1860 2864 1912 2916
rect 32128 2941 32137 2975
rect 32137 2941 32171 2975
rect 32171 2941 32180 2975
rect 32128 2932 32180 2941
rect 40132 3000 40184 3052
rect 43352 3043 43404 3052
rect 43352 3009 43361 3043
rect 43361 3009 43395 3043
rect 43395 3009 43404 3043
rect 43352 3000 43404 3009
rect 52828 3068 52880 3120
rect 46388 3000 46440 3052
rect 47768 3043 47820 3052
rect 47768 3009 47777 3043
rect 47777 3009 47811 3043
rect 47811 3009 47820 3043
rect 47768 3000 47820 3009
rect 35624 2932 35676 2984
rect 39672 2932 39724 2984
rect 39856 2975 39908 2984
rect 39856 2941 39865 2975
rect 39865 2941 39899 2975
rect 39899 2941 39908 2975
rect 43168 2975 43220 2984
rect 39856 2932 39908 2941
rect 43168 2941 43177 2975
rect 43177 2941 43211 2975
rect 43211 2941 43220 2975
rect 43168 2932 43220 2941
rect 43628 2932 43680 2984
rect 47584 2975 47636 2984
rect 47584 2941 47593 2975
rect 47593 2941 47627 2975
rect 47627 2941 47636 2975
rect 47584 2932 47636 2941
rect 1124 2796 1176 2848
rect 2780 2796 2832 2848
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 28356 2796 28408 2848
rect 29092 2796 29144 2848
rect 31576 2839 31628 2848
rect 31576 2805 31585 2839
rect 31585 2805 31619 2839
rect 31619 2805 31628 2839
rect 31576 2796 31628 2805
rect 32864 2796 32916 2848
rect 35440 2796 35492 2848
rect 35532 2796 35584 2848
rect 37096 2796 37148 2848
rect 39488 2796 39540 2848
rect 40224 2839 40276 2848
rect 40224 2805 40233 2839
rect 40233 2805 40267 2839
rect 40267 2805 40276 2839
rect 40224 2796 40276 2805
rect 50620 3043 50672 3052
rect 50620 3009 50629 3043
rect 50629 3009 50663 3043
rect 50663 3009 50672 3043
rect 50620 3000 50672 3009
rect 52368 3000 52420 3052
rect 53288 3145 53297 3179
rect 53297 3145 53331 3179
rect 53331 3145 53340 3179
rect 53288 3136 53340 3145
rect 54944 3179 54996 3188
rect 54944 3145 54953 3179
rect 54953 3145 54987 3179
rect 54987 3145 54996 3179
rect 54944 3136 54996 3145
rect 53012 3000 53064 3052
rect 56600 3000 56652 3052
rect 57980 3136 58032 3188
rect 62396 3136 62448 3188
rect 66352 3179 66404 3188
rect 66352 3145 66361 3179
rect 66361 3145 66395 3179
rect 66395 3145 66404 3179
rect 66352 3136 66404 3145
rect 68376 3179 68428 3188
rect 68376 3145 68385 3179
rect 68385 3145 68419 3179
rect 68419 3145 68428 3179
rect 68376 3136 68428 3145
rect 83556 3136 83608 3188
rect 112628 3136 112680 3188
rect 56968 3111 57020 3120
rect 56968 3077 56977 3111
rect 56977 3077 57011 3111
rect 57011 3077 57020 3111
rect 56968 3068 57020 3077
rect 61844 3068 61896 3120
rect 56784 3043 56836 3052
rect 56784 3009 56793 3043
rect 56793 3009 56827 3043
rect 56827 3009 56836 3043
rect 56784 3000 56836 3009
rect 57152 3000 57204 3052
rect 59544 3000 59596 3052
rect 61936 3000 61988 3052
rect 79140 3068 79192 3120
rect 66260 3043 66312 3052
rect 66260 3009 66269 3043
rect 66269 3009 66303 3043
rect 66303 3009 66312 3043
rect 66260 3000 66312 3009
rect 68192 3043 68244 3052
rect 68192 3009 68201 3043
rect 68201 3009 68235 3043
rect 68235 3009 68244 3043
rect 68192 3000 68244 3009
rect 73620 3043 73672 3052
rect 54852 2932 54904 2984
rect 57336 2932 57388 2984
rect 46204 2796 46256 2848
rect 46296 2796 46348 2848
rect 57428 2864 57480 2916
rect 50712 2796 50764 2848
rect 51908 2796 51960 2848
rect 68652 2932 68704 2984
rect 70768 2975 70820 2984
rect 70768 2941 70777 2975
rect 70777 2941 70811 2975
rect 70811 2941 70820 2975
rect 70768 2932 70820 2941
rect 73620 3009 73629 3043
rect 73629 3009 73663 3043
rect 73663 3009 73672 3043
rect 73620 3000 73672 3009
rect 73712 3000 73764 3052
rect 76288 3000 76340 3052
rect 76748 3000 76800 3052
rect 83648 3043 83700 3052
rect 79968 2975 80020 2984
rect 79968 2941 79977 2975
rect 79977 2941 80011 2975
rect 80011 2941 80020 2975
rect 79968 2932 80020 2941
rect 83648 3009 83657 3043
rect 83657 3009 83691 3043
rect 83691 3009 83700 3043
rect 83648 3000 83700 3009
rect 85948 3000 86000 3052
rect 86868 3043 86920 3052
rect 86868 3009 86877 3043
rect 86877 3009 86911 3043
rect 86911 3009 86920 3043
rect 86868 3000 86920 3009
rect 88156 3000 88208 3052
rect 89628 3068 89680 3120
rect 93860 3068 93912 3120
rect 94964 3068 95016 3120
rect 95056 3068 95108 3120
rect 89352 3043 89404 3052
rect 89352 3009 89361 3043
rect 89361 3009 89395 3043
rect 89395 3009 89404 3043
rect 89352 3000 89404 3009
rect 91192 3043 91244 3052
rect 91192 3009 91201 3043
rect 91201 3009 91235 3043
rect 91235 3009 91244 3043
rect 91192 3000 91244 3009
rect 92020 3043 92072 3052
rect 92020 3009 92029 3043
rect 92029 3009 92063 3043
rect 92063 3009 92072 3043
rect 92020 3000 92072 3009
rect 94044 3000 94096 3052
rect 96896 3000 96948 3052
rect 99564 3043 99616 3052
rect 99564 3009 99573 3043
rect 99573 3009 99607 3043
rect 99607 3009 99616 3043
rect 99564 3000 99616 3009
rect 100392 3000 100444 3052
rect 104256 3043 104308 3052
rect 104256 3009 104265 3043
rect 104265 3009 104299 3043
rect 104299 3009 104308 3043
rect 104256 3000 104308 3009
rect 104992 3000 105044 3052
rect 107292 3043 107344 3052
rect 107292 3009 107301 3043
rect 107301 3009 107335 3043
rect 107335 3009 107344 3043
rect 107292 3000 107344 3009
rect 108304 3000 108356 3052
rect 57612 2864 57664 2916
rect 73988 2864 74040 2916
rect 62028 2796 62080 2848
rect 62120 2796 62172 2848
rect 65156 2796 65208 2848
rect 74632 2796 74684 2848
rect 74724 2796 74776 2848
rect 76380 2839 76432 2848
rect 76380 2805 76389 2839
rect 76389 2805 76423 2839
rect 76423 2805 76432 2839
rect 76380 2796 76432 2805
rect 77116 2796 77168 2848
rect 81900 2796 81952 2848
rect 98000 2932 98052 2984
rect 90640 2864 90692 2916
rect 91744 2864 91796 2916
rect 87696 2796 87748 2848
rect 87972 2796 88024 2848
rect 89352 2796 89404 2848
rect 90272 2839 90324 2848
rect 90272 2805 90281 2839
rect 90281 2805 90315 2839
rect 90315 2805 90324 2839
rect 90272 2796 90324 2805
rect 92112 2839 92164 2848
rect 92112 2805 92121 2839
rect 92121 2805 92155 2839
rect 92155 2805 92164 2839
rect 92112 2796 92164 2805
rect 96988 2864 97040 2916
rect 105176 2864 105228 2916
rect 96252 2796 96304 2848
rect 99472 2796 99524 2848
rect 100944 2796 100996 2848
rect 103520 2796 103572 2848
rect 105084 2796 105136 2848
rect 109776 2864 109828 2916
rect 115572 3136 115624 3188
rect 111432 3000 111484 3052
rect 112260 3000 112312 3052
rect 114836 3043 114888 3052
rect 114836 3009 114845 3043
rect 114845 3009 114879 3043
rect 114879 3009 114888 3043
rect 114836 3000 114888 3009
rect 117964 3043 118016 3052
rect 117964 3009 117973 3043
rect 117973 3009 118007 3043
rect 118007 3009 118016 3043
rect 117964 3000 118016 3009
rect 110972 2932 111024 2984
rect 109960 2796 110012 2848
rect 112168 2796 112220 2848
rect 114744 2796 114796 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 22376 2635 22428 2644
rect 22376 2601 22385 2635
rect 22385 2601 22419 2635
rect 22419 2601 22428 2635
rect 22376 2592 22428 2601
rect 23480 2592 23532 2644
rect 28632 2592 28684 2644
rect 30840 2592 30892 2644
rect 37832 2592 37884 2644
rect 2412 2499 2464 2508
rect 2412 2465 2421 2499
rect 2421 2465 2455 2499
rect 2455 2465 2464 2499
rect 2412 2456 2464 2465
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 4344 2388 4396 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5908 2388 5960 2440
rect 9128 2388 9180 2440
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10784 2388 10836 2440
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 33140 2524 33192 2576
rect 43168 2592 43220 2644
rect 43260 2592 43312 2644
rect 15568 2388 15620 2440
rect 7564 2320 7616 2372
rect 12348 2320 12400 2372
rect 34060 2456 34112 2508
rect 17132 2388 17184 2440
rect 18696 2431 18748 2440
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 19432 2388 19484 2440
rect 20352 2388 20404 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 23480 2388 23532 2440
rect 23572 2388 23624 2440
rect 24400 2431 24452 2440
rect 24400 2397 24409 2431
rect 24409 2397 24443 2431
rect 24443 2397 24452 2431
rect 24400 2388 24452 2397
rect 25136 2388 25188 2440
rect 26700 2388 26752 2440
rect 27528 2388 27580 2440
rect 28632 2431 28684 2440
rect 3516 2252 3568 2304
rect 5172 2252 5224 2304
rect 7840 2295 7892 2304
rect 7840 2261 7849 2295
rect 7849 2261 7883 2295
rect 7883 2261 7892 2295
rect 7840 2252 7892 2261
rect 9956 2252 10008 2304
rect 13176 2252 13228 2304
rect 14740 2252 14792 2304
rect 26884 2320 26936 2372
rect 28632 2397 28641 2431
rect 28641 2397 28675 2431
rect 28675 2397 28684 2431
rect 28632 2388 28684 2397
rect 30748 2388 30800 2440
rect 31668 2431 31720 2440
rect 31668 2397 31677 2431
rect 31677 2397 31711 2431
rect 31711 2397 31720 2431
rect 31668 2388 31720 2397
rect 32864 2431 32916 2440
rect 32864 2397 32873 2431
rect 32873 2397 32907 2431
rect 32907 2397 32916 2431
rect 32864 2388 32916 2397
rect 45468 2592 45520 2644
rect 52276 2592 52328 2644
rect 52460 2592 52512 2644
rect 53196 2592 53248 2644
rect 85396 2635 85448 2644
rect 34244 2456 34296 2508
rect 39856 2456 39908 2508
rect 34980 2431 35032 2440
rect 17960 2252 18012 2304
rect 19432 2252 19484 2304
rect 22744 2252 22796 2304
rect 24308 2252 24360 2304
rect 34980 2397 34989 2431
rect 34989 2397 35023 2431
rect 35023 2397 35032 2431
rect 34980 2388 35032 2397
rect 30656 2295 30708 2304
rect 30656 2261 30665 2295
rect 30665 2261 30699 2295
rect 30699 2261 30708 2295
rect 30656 2252 30708 2261
rect 32312 2252 32364 2304
rect 33232 2320 33284 2372
rect 35072 2320 35124 2372
rect 36544 2363 36596 2372
rect 36544 2329 36553 2363
rect 36553 2329 36587 2363
rect 36587 2329 36596 2363
rect 36544 2320 36596 2329
rect 38752 2388 38804 2440
rect 43260 2456 43312 2508
rect 61752 2524 61804 2576
rect 61936 2567 61988 2576
rect 61936 2533 61945 2567
rect 61945 2533 61979 2567
rect 61979 2533 61988 2567
rect 61936 2524 61988 2533
rect 62028 2524 62080 2576
rect 40684 2431 40736 2440
rect 40684 2397 40693 2431
rect 40693 2397 40727 2431
rect 40727 2397 40736 2431
rect 40684 2388 40736 2397
rect 41144 2388 41196 2440
rect 42708 2388 42760 2440
rect 43444 2388 43496 2440
rect 44088 2388 44140 2440
rect 45100 2388 45152 2440
rect 45928 2388 45980 2440
rect 47492 2388 47544 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 48320 2388 48372 2440
rect 49884 2388 49936 2440
rect 62672 2456 62724 2508
rect 64052 2524 64104 2576
rect 65800 2524 65852 2576
rect 66260 2524 66312 2576
rect 67548 2524 67600 2576
rect 33692 2295 33744 2304
rect 33692 2261 33701 2295
rect 33701 2261 33735 2295
rect 33735 2261 33744 2295
rect 33692 2252 33744 2261
rect 36360 2252 36412 2304
rect 38384 2295 38436 2304
rect 38384 2261 38393 2295
rect 38393 2261 38427 2295
rect 38427 2261 38436 2295
rect 38384 2252 38436 2261
rect 39212 2295 39264 2304
rect 39212 2261 39221 2295
rect 39221 2261 39255 2295
rect 39255 2261 39264 2295
rect 39212 2252 39264 2261
rect 40040 2252 40092 2304
rect 40408 2252 40460 2304
rect 44088 2252 44140 2304
rect 52276 2388 52328 2440
rect 53012 2388 53064 2440
rect 53104 2388 53156 2440
rect 54760 2431 54812 2440
rect 54760 2397 54769 2431
rect 54769 2397 54803 2431
rect 54803 2397 54812 2431
rect 54760 2388 54812 2397
rect 55496 2388 55548 2440
rect 56600 2431 56652 2440
rect 53196 2320 53248 2372
rect 46848 2295 46900 2304
rect 46848 2261 46857 2295
rect 46857 2261 46891 2295
rect 46891 2261 46900 2295
rect 46848 2252 46900 2261
rect 53012 2252 53064 2304
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 57888 2388 57940 2440
rect 60372 2388 60424 2440
rect 66812 2499 66864 2508
rect 66812 2465 66821 2499
rect 66821 2465 66855 2499
rect 66855 2465 66864 2499
rect 66812 2456 66864 2465
rect 68836 2499 68888 2508
rect 62120 2320 62172 2372
rect 62764 2320 62816 2372
rect 64328 2388 64380 2440
rect 65800 2431 65852 2440
rect 59820 2295 59872 2304
rect 59820 2261 59829 2295
rect 59829 2261 59863 2295
rect 59863 2261 59872 2295
rect 59820 2252 59872 2261
rect 65800 2397 65809 2431
rect 65809 2397 65843 2431
rect 65843 2397 65852 2431
rect 65800 2388 65852 2397
rect 66720 2388 66772 2440
rect 68836 2465 68845 2499
rect 68845 2465 68879 2499
rect 68879 2465 68888 2499
rect 68836 2456 68888 2465
rect 68652 2431 68704 2440
rect 68652 2397 68661 2431
rect 68661 2397 68695 2431
rect 68695 2397 68704 2431
rect 68652 2388 68704 2397
rect 73712 2567 73764 2576
rect 70032 2456 70084 2508
rect 73712 2533 73721 2567
rect 73721 2533 73755 2567
rect 73755 2533 73764 2567
rect 73712 2524 73764 2533
rect 70124 2431 70176 2440
rect 65708 2252 65760 2304
rect 70124 2397 70133 2431
rect 70133 2397 70167 2431
rect 70167 2397 70176 2431
rect 70124 2388 70176 2397
rect 71504 2388 71556 2440
rect 72332 2388 72384 2440
rect 70768 2320 70820 2372
rect 74540 2499 74592 2508
rect 74540 2465 74549 2499
rect 74549 2465 74583 2499
rect 74583 2465 74592 2499
rect 74540 2456 74592 2465
rect 76380 2456 76432 2508
rect 79048 2524 79100 2576
rect 79968 2524 80020 2576
rect 81992 2456 82044 2508
rect 78680 2388 78732 2440
rect 79508 2388 79560 2440
rect 81348 2388 81400 2440
rect 85396 2601 85405 2635
rect 85405 2601 85439 2635
rect 85439 2601 85448 2635
rect 85396 2592 85448 2601
rect 88156 2635 88208 2644
rect 88156 2601 88165 2635
rect 88165 2601 88199 2635
rect 88199 2601 88208 2635
rect 88156 2592 88208 2601
rect 89444 2635 89496 2644
rect 89444 2601 89453 2635
rect 89453 2601 89487 2635
rect 89487 2601 89496 2635
rect 89444 2592 89496 2601
rect 91836 2592 91888 2644
rect 91928 2592 91980 2644
rect 96896 2635 96948 2644
rect 96896 2601 96905 2635
rect 96905 2601 96939 2635
rect 96939 2601 96948 2635
rect 96896 2592 96948 2601
rect 104992 2592 105044 2644
rect 108304 2635 108356 2644
rect 108304 2601 108313 2635
rect 108313 2601 108347 2635
rect 108347 2601 108356 2635
rect 108304 2592 108356 2601
rect 112260 2592 112312 2644
rect 79048 2320 79100 2372
rect 76104 2295 76156 2304
rect 76104 2261 76113 2295
rect 76113 2261 76147 2295
rect 76147 2261 76156 2295
rect 76104 2252 76156 2261
rect 79140 2252 79192 2304
rect 83556 2388 83608 2440
rect 84292 2388 84344 2440
rect 98092 2524 98144 2576
rect 84844 2456 84896 2508
rect 90456 2456 90508 2508
rect 87972 2431 88024 2440
rect 87972 2397 87981 2431
rect 87981 2397 88015 2431
rect 88015 2397 88024 2431
rect 87972 2388 88024 2397
rect 88156 2388 88208 2440
rect 89628 2431 89680 2440
rect 89628 2397 89637 2431
rect 89637 2397 89671 2431
rect 89671 2397 89680 2431
rect 89628 2388 89680 2397
rect 90548 2431 90600 2440
rect 90548 2397 90557 2431
rect 90557 2397 90591 2431
rect 90591 2397 90600 2431
rect 90548 2388 90600 2397
rect 90640 2431 90692 2440
rect 90640 2397 90649 2431
rect 90649 2397 90683 2431
rect 90683 2397 90692 2431
rect 91652 2456 91704 2508
rect 93952 2456 94004 2508
rect 100300 2524 100352 2576
rect 99012 2456 99064 2508
rect 102324 2456 102376 2508
rect 109960 2499 110012 2508
rect 109960 2465 109969 2499
rect 109969 2465 110003 2499
rect 110003 2465 110012 2499
rect 109960 2456 110012 2465
rect 90640 2388 90692 2397
rect 86776 2295 86828 2304
rect 86776 2261 86785 2295
rect 86785 2261 86819 2295
rect 86819 2261 86828 2295
rect 86776 2252 86828 2261
rect 89444 2320 89496 2372
rect 92388 2431 92440 2440
rect 92388 2397 92397 2431
rect 92397 2397 92431 2431
rect 92431 2397 92440 2431
rect 92388 2388 92440 2397
rect 93400 2388 93452 2440
rect 95516 2388 95568 2440
rect 96712 2431 96764 2440
rect 92020 2252 92072 2304
rect 92388 2252 92440 2304
rect 96712 2397 96721 2431
rect 96721 2397 96755 2431
rect 96755 2397 96764 2431
rect 96712 2388 96764 2397
rect 97908 2388 97960 2440
rect 100944 2431 100996 2440
rect 100944 2397 100953 2431
rect 100953 2397 100987 2431
rect 100987 2397 100996 2431
rect 100944 2388 100996 2397
rect 100392 2252 100444 2304
rect 102784 2431 102836 2440
rect 102784 2397 102793 2431
rect 102793 2397 102827 2431
rect 102827 2397 102836 2431
rect 102784 2388 102836 2397
rect 104900 2431 104952 2440
rect 104900 2397 104934 2431
rect 104934 2397 104952 2431
rect 104900 2388 104952 2397
rect 107568 2431 107620 2440
rect 107568 2397 107577 2431
rect 107577 2397 107611 2431
rect 107611 2397 107620 2431
rect 107568 2388 107620 2397
rect 109776 2431 109828 2440
rect 101220 2295 101272 2304
rect 101220 2261 101229 2295
rect 101229 2261 101263 2295
rect 101263 2261 101272 2295
rect 101220 2252 101272 2261
rect 102692 2252 102744 2304
rect 107476 2252 107528 2304
rect 109776 2397 109785 2431
rect 109785 2397 109819 2431
rect 109819 2397 109828 2431
rect 109776 2388 109828 2397
rect 109868 2388 109920 2440
rect 112076 2388 112128 2440
rect 110696 2320 110748 2372
rect 112352 2524 112404 2576
rect 112812 2388 112864 2440
rect 114560 2431 114612 2440
rect 114560 2397 114569 2431
rect 114569 2397 114603 2431
rect 114603 2397 114612 2431
rect 114560 2388 114612 2397
rect 115480 2388 115532 2440
rect 115848 2431 115900 2440
rect 115848 2397 115857 2431
rect 115857 2397 115891 2431
rect 115891 2397 115900 2431
rect 115848 2388 115900 2397
rect 117136 2431 117188 2440
rect 117136 2397 117145 2431
rect 117145 2397 117179 2431
rect 117179 2397 117188 2431
rect 117136 2388 117188 2397
rect 117228 2388 117280 2440
rect 117412 2320 117464 2372
rect 112812 2295 112864 2304
rect 112812 2261 112821 2295
rect 112821 2261 112855 2295
rect 112855 2261 112864 2295
rect 112812 2252 112864 2261
rect 113916 2252 113968 2304
rect 116308 2252 116360 2304
rect 117872 2252 117924 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 81014 2150 81066 2202
rect 81078 2150 81130 2202
rect 81142 2150 81194 2202
rect 81206 2150 81258 2202
rect 81270 2150 81322 2202
rect 111734 2150 111786 2202
rect 111798 2150 111850 2202
rect 111862 2150 111914 2202
rect 111926 2150 111978 2202
rect 111990 2150 112042 2202
rect 26884 2048 26936 2100
rect 32128 2048 32180 2100
rect 35072 2048 35124 2100
rect 39212 2048 39264 2100
rect 44088 2048 44140 2100
rect 47768 2048 47820 2100
rect 59820 2048 59872 2100
rect 107568 2048 107620 2100
rect 7840 1980 7892 2032
rect 34980 1980 35032 2032
rect 46848 1980 46900 2032
rect 54852 1980 54904 2032
rect 76104 1980 76156 2032
rect 114560 1980 114612 2032
rect 38384 1912 38436 1964
rect 46480 1912 46532 1964
rect 81992 1912 82044 1964
rect 84844 1912 84896 1964
rect 86776 1912 86828 1964
rect 117228 1912 117280 1964
rect 85396 1844 85448 1896
rect 117136 1844 117188 1896
rect 90456 1776 90508 1828
rect 96712 1776 96764 1828
rect 99380 1776 99432 1828
rect 115848 1776 115900 1828
rect 30656 1708 30708 1760
rect 102784 1708 102836 1760
rect 36544 1640 36596 1692
rect 99564 1640 99616 1692
rect 79140 1572 79192 1624
rect 114836 1572 114888 1624
rect 33692 1504 33744 1556
rect 101220 1504 101272 1556
rect 74632 1436 74684 1488
rect 112812 1436 112864 1488
rect 69112 1368 69164 1420
rect 70124 1368 70176 1420
rect 86684 1368 86736 1420
rect 88156 1368 88208 1420
rect 88340 1368 88392 1420
rect 89628 1368 89680 1420
<< metal2 >>
rect 2042 39200 2098 40000
rect 6090 39200 6146 40000
rect 10230 39200 10286 40000
rect 14370 39200 14426 40000
rect 18510 39200 18566 40000
rect 22650 39200 22706 40000
rect 26790 39200 26846 40000
rect 30930 39200 30986 40000
rect 35070 39200 35126 40000
rect 35176 39222 35388 39250
rect 1582 37496 1638 37505
rect 2056 37466 2084 39200
rect 2778 39128 2834 39137
rect 2778 39063 2834 39072
rect 1582 37431 1584 37440
rect 1636 37431 1638 37440
rect 2044 37460 2096 37466
rect 1584 37402 1636 37408
rect 2044 37402 2096 37408
rect 2792 36922 2820 39063
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 10244 37262 10272 39200
rect 14384 37466 14412 39200
rect 22664 37466 22692 39200
rect 26804 37466 26832 39200
rect 30944 37466 30972 39200
rect 35084 39114 35112 39200
rect 35176 39114 35204 39222
rect 35084 39086 35204 39114
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 37466 35388 39222
rect 39210 39200 39266 40000
rect 43350 39200 43406 40000
rect 47490 39200 47546 40000
rect 51630 39200 51686 40000
rect 55770 39200 55826 40000
rect 59910 39200 59966 40000
rect 64050 39200 64106 40000
rect 68190 39200 68246 40000
rect 72330 39200 72386 40000
rect 76470 39200 76526 40000
rect 80610 39200 80666 40000
rect 84750 39200 84806 40000
rect 88890 39200 88946 40000
rect 93030 39200 93086 40000
rect 97170 39200 97226 40000
rect 101310 39200 101366 40000
rect 105450 39200 105506 40000
rect 109590 39200 109646 40000
rect 113730 39200 113786 40000
rect 117226 39264 117282 39273
rect 14372 37460 14424 37466
rect 14372 37402 14424 37408
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 26792 37460 26844 37466
rect 26792 37402 26844 37408
rect 30932 37460 30984 37466
rect 30932 37402 30984 37408
rect 35348 37460 35400 37466
rect 35348 37402 35400 37408
rect 39224 37262 39252 39200
rect 10232 37256 10284 37262
rect 10232 37198 10284 37204
rect 39212 37256 39264 37262
rect 39212 37198 39264 37204
rect 40500 37188 40552 37194
rect 40500 37130 40552 37136
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 2780 36916 2832 36922
rect 2780 36858 2832 36864
rect 40512 36854 40540 37130
rect 47504 37126 47532 39200
rect 50896 37324 50948 37330
rect 50896 37266 50948 37272
rect 47584 37256 47636 37262
rect 47584 37198 47636 37204
rect 47492 37120 47544 37126
rect 47492 37062 47544 37068
rect 45560 36916 45612 36922
rect 45560 36858 45612 36864
rect 40500 36848 40552 36854
rect 40500 36790 40552 36796
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 1492 36168 1544 36174
rect 1492 36110 1544 36116
rect 1504 35873 1532 36110
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 1490 35864 1546 35873
rect 19574 35867 19882 35876
rect 1490 35799 1546 35808
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 26042 1440 34546
rect 1584 34400 1636 34406
rect 1584 34342 1636 34348
rect 1596 34241 1624 34342
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 1582 34232 1638 34241
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 1582 34167 1638 34176
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25809 1440 25842
rect 1398 25800 1454 25809
rect 1398 25735 1454 25744
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22545 1440 22578
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19145 1440 19314
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 17513 1440 17614
rect 1398 17504 1454 17513
rect 1398 17439 1454 17448
rect 1504 17082 1532 32846
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1596 32473 1624 32710
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 1582 32464 1638 32473
rect 1582 32399 1638 32408
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 1596 29209 1624 29446
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1768 26036 1820 26042
rect 1768 25978 1820 25984
rect 1676 25832 1728 25838
rect 1676 25774 1728 25780
rect 1582 24168 1638 24177
rect 1582 24103 1638 24112
rect 1596 24070 1624 24103
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1688 20398 1716 25774
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19446 1716 19654
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 1780 19334 1808 25978
rect 1860 24200 1912 24206
rect 1860 24142 1912 24148
rect 1320 17054 1532 17082
rect 1596 19306 1808 19334
rect 1320 14550 1348 17054
rect 1596 14634 1624 19306
rect 1872 17626 1900 24142
rect 1412 14606 1624 14634
rect 1688 17598 1900 17626
rect 1308 14544 1360 14550
rect 1308 14486 1360 14492
rect 1412 4146 1440 14606
rect 1492 14544 1544 14550
rect 1492 14486 1544 14492
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 388 3392 440 3398
rect 388 3334 440 3340
rect 400 800 428 3334
rect 1412 3194 1440 3470
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1504 3126 1532 14486
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 9217 1624 9318
rect 1582 9208 1638 9217
rect 1582 9143 1638 9152
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7585 1624 7822
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 1688 3602 1716 17598
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1780 5030 1808 17478
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1872 14249 1900 14282
rect 1952 14272 2004 14278
rect 1858 14240 1914 14249
rect 1952 14214 2004 14220
rect 1858 14175 1914 14184
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1872 10849 1900 11018
rect 1858 10840 1914 10849
rect 1858 10775 1914 10784
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1492 3120 1544 3126
rect 1492 3062 1544 3068
rect 1872 2922 1900 10678
rect 1964 5098 1992 14214
rect 2056 10742 2084 29582
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 45572 16574 45600 36858
rect 45572 16546 45692 16574
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 39672 12096 39724 12102
rect 39672 12038 39724 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 2044 10736 2096 10742
rect 2044 10678 2096 10684
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 7576 5302 7604 11018
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 22112 8430 22140 9522
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2424 3534 2452 4558
rect 9876 4554 9904 5510
rect 10060 5370 10088 5646
rect 10336 5370 10364 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 10244 4486 10272 5170
rect 17144 4622 17172 5510
rect 17236 5370 17264 5646
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18432 4826 18460 5170
rect 20824 5030 20852 5306
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4146 10272 4422
rect 18432 4146 18460 4762
rect 21376 4622 21404 4966
rect 22204 4826 22232 5170
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 2608 3534 2636 4082
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1124 2848 1176 2854
rect 1124 2790 1176 2796
rect 1136 800 1164 2790
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 921 1440 2382
rect 1398 912 1454 921
rect 1398 847 1454 856
rect 1964 800 1992 3402
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3058 2268 3334
rect 2424 3058 2452 3470
rect 2884 3058 2912 3674
rect 10152 3534 10180 3878
rect 19996 3534 20024 3878
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 2424 2514 2452 2994
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2792 800 2820 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5276 2446 5304 2994
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 800 3556 2246
rect 4356 800 4384 2382
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5920 800 5948 2382
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7576 800 7604 2314
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 7852 2038 7880 2246
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 8312 800 8340 2926
rect 10060 2446 10088 3334
rect 19444 2446 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 9140 800 9168 2382
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 800 9996 2246
rect 10796 800 10824 2382
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12360 800 12388 2314
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13188 800 13216 2246
rect 13924 800 13952 2382
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 800 14780 2246
rect 15580 800 15608 2382
rect 17144 800 17172 2382
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 800 18000 2246
rect 18708 800 18736 2382
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 1170 19472 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1142 19564 1170
rect 19536 800 19564 1142
rect 20364 800 20392 2382
rect 21928 800 21956 2994
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22020 2446 22048 2790
rect 22388 2650 22416 8434
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 39684 5370 39712 12038
rect 39672 5364 39724 5370
rect 39672 5306 39724 5312
rect 39856 5364 39908 5370
rect 39856 5306 39908 5312
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 39580 5228 39632 5234
rect 39580 5170 39632 5176
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22756 4078 22784 4762
rect 28644 4486 28672 5170
rect 29736 5024 29788 5030
rect 29736 4966 29788 4972
rect 38660 5024 38712 5030
rect 38660 4966 38712 4972
rect 29748 4622 29776 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 38568 4820 38620 4826
rect 38568 4762 38620 4768
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28632 4480 28684 4486
rect 28632 4422 28684 4428
rect 28184 4078 28212 4422
rect 38580 4078 38608 4762
rect 38672 4146 38700 4966
rect 39592 4282 39620 5170
rect 39868 5166 39896 5306
rect 39856 5160 39908 5166
rect 39856 5102 39908 5108
rect 38752 4276 38804 4282
rect 38752 4218 38804 4224
rect 39580 4276 39632 4282
rect 39580 4218 39632 4224
rect 38660 4140 38712 4146
rect 38660 4082 38712 4088
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 28172 4072 28224 4078
rect 28172 4014 28224 4020
rect 38568 4072 38620 4078
rect 38568 4014 38620 4020
rect 35348 4004 35400 4010
rect 35348 3946 35400 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 23768 3534 23796 3878
rect 28552 3534 28580 3878
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23492 2446 23520 2586
rect 24412 2446 24440 3334
rect 28460 3058 28488 3334
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22756 800 22784 2246
rect 23584 800 23612 2382
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 24320 800 24348 2246
rect 25148 800 25176 2382
rect 26712 800 26740 2382
rect 26884 2372 26936 2378
rect 26884 2314 26936 2320
rect 26896 2106 26924 2314
rect 26884 2100 26936 2106
rect 26884 2042 26936 2048
rect 27540 800 27568 2382
rect 28368 800 28396 2790
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28644 2446 28672 2586
rect 28632 2440 28684 2446
rect 28632 2382 28684 2388
rect 29104 800 29132 2790
rect 30852 2650 30880 2994
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 30656 2304 30708 2310
rect 30656 2246 30708 2252
rect 30668 1766 30696 2246
rect 30656 1760 30708 1766
rect 30656 1702 30708 1708
rect 30760 800 30788 2382
rect 31588 800 31616 2790
rect 31680 2446 31708 3878
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35360 3670 35388 3946
rect 35348 3664 35400 3670
rect 35348 3606 35400 3612
rect 38384 3664 38436 3670
rect 38764 3618 38792 4218
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 42892 3936 42944 3942
rect 42892 3878 42944 3884
rect 38384 3606 38436 3612
rect 37832 3460 37884 3466
rect 37832 3402 37884 3408
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 34704 3052 34756 3058
rect 34704 2994 34756 3000
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 32140 2106 32168 2926
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32876 2446 32904 2790
rect 33060 2666 33088 2994
rect 33060 2638 33272 2666
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 32128 2100 32180 2106
rect 32128 2042 32180 2048
rect 32324 800 32352 2246
rect 33152 800 33180 2518
rect 33244 2378 33272 2638
rect 34072 2514 34284 2530
rect 34060 2508 34296 2514
rect 34112 2502 34244 2508
rect 34060 2450 34112 2456
rect 34244 2450 34296 2456
rect 33232 2372 33284 2378
rect 33232 2314 33284 2320
rect 33692 2304 33744 2310
rect 33692 2246 33744 2252
rect 33704 1562 33732 2246
rect 33692 1556 33744 1562
rect 33692 1498 33744 1504
rect 34716 800 34744 2994
rect 35624 2984 35676 2990
rect 35452 2932 35624 2938
rect 35452 2926 35676 2932
rect 35452 2910 35664 2926
rect 35452 2854 35480 2910
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 37096 2848 37148 2854
rect 37096 2790 37148 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 34992 2038 35020 2382
rect 35072 2372 35124 2378
rect 35072 2314 35124 2320
rect 35084 2106 35112 2314
rect 35072 2100 35124 2106
rect 35072 2042 35124 2048
rect 34980 2032 35032 2038
rect 34980 1974 35032 1980
rect 35544 800 35572 2790
rect 36544 2372 36596 2378
rect 36544 2314 36596 2320
rect 36360 2304 36412 2310
rect 36360 2246 36412 2252
rect 36372 800 36400 2246
rect 36556 1698 36584 2314
rect 36544 1692 36596 1698
rect 36544 1634 36596 1640
rect 37108 800 37136 2790
rect 37844 2650 37872 3402
rect 38396 3346 38424 3606
rect 38488 3590 38792 3618
rect 38488 3534 38516 3590
rect 42904 3534 42932 3878
rect 45480 3670 45508 4014
rect 45664 3670 45692 16546
rect 47596 3670 47624 37198
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50908 5370 50936 37266
rect 51644 37262 51672 39200
rect 51632 37256 51684 37262
rect 51632 37198 51684 37204
rect 54944 37256 54996 37262
rect 54944 37198 54996 37204
rect 54116 23520 54168 23526
rect 54116 23462 54168 23468
rect 52736 22432 52788 22438
rect 52736 22374 52788 22380
rect 49884 5364 49936 5370
rect 49884 5306 49936 5312
rect 49976 5364 50028 5370
rect 50068 5364 50120 5370
rect 50028 5324 50068 5352
rect 49976 5306 50028 5312
rect 50068 5306 50120 5312
rect 50896 5364 50948 5370
rect 50896 5306 50948 5312
rect 49332 5228 49384 5234
rect 49332 5170 49384 5176
rect 48596 5160 48648 5166
rect 48596 5102 48648 5108
rect 48608 5030 48636 5102
rect 48596 5024 48648 5030
rect 48596 4966 48648 4972
rect 48608 4826 48636 4966
rect 49344 4826 49372 5170
rect 49896 5166 49924 5306
rect 49884 5160 49936 5166
rect 49884 5102 49936 5108
rect 48596 4820 48648 4826
rect 48596 4762 48648 4768
rect 49332 4820 49384 4826
rect 49332 4762 49384 4768
rect 49988 4690 50016 5306
rect 50988 5160 51040 5166
rect 50988 5102 51040 5108
rect 50068 5024 50120 5030
rect 50068 4966 50120 4972
rect 49976 4684 50028 4690
rect 49976 4626 50028 4632
rect 50080 4622 50108 4966
rect 51000 4690 51028 5102
rect 50988 4684 51040 4690
rect 50988 4626 51040 4632
rect 50068 4616 50120 4622
rect 50068 4558 50120 4564
rect 50620 4616 50672 4622
rect 50620 4558 50672 4564
rect 50160 4480 50212 4486
rect 50160 4422 50212 4428
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47688 3670 47716 3878
rect 45468 3664 45520 3670
rect 45468 3606 45520 3612
rect 45652 3664 45704 3670
rect 45652 3606 45704 3612
rect 47584 3664 47636 3670
rect 47584 3606 47636 3612
rect 47676 3664 47728 3670
rect 47676 3606 47728 3612
rect 50172 3534 50200 4422
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50632 4078 50660 4558
rect 50620 4072 50672 4078
rect 50620 4014 50672 4020
rect 52460 3936 52512 3942
rect 52460 3878 52512 3884
rect 52472 3670 52500 3878
rect 52460 3664 52512 3670
rect 52460 3606 52512 3612
rect 52748 3602 52776 22374
rect 53564 5228 53616 5234
rect 53564 5170 53616 5176
rect 53576 4622 53604 5170
rect 53564 4616 53616 4622
rect 53564 4558 53616 4564
rect 53576 4282 53604 4558
rect 53564 4276 53616 4282
rect 53564 4218 53616 4224
rect 54128 3602 54156 23462
rect 52736 3596 52788 3602
rect 52736 3538 52788 3544
rect 54116 3596 54168 3602
rect 54116 3538 54168 3544
rect 38476 3528 38528 3534
rect 38476 3470 38528 3476
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 46480 3528 46532 3534
rect 46480 3470 46532 3476
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 52460 3528 52512 3534
rect 52460 3470 52512 3476
rect 52828 3528 52880 3534
rect 52828 3470 52880 3476
rect 38580 3346 38608 3470
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 38396 3318 38608 3346
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 39672 2984 39724 2990
rect 39670 2952 39672 2961
rect 39856 2984 39908 2990
rect 39724 2952 39726 2961
rect 39856 2926 39908 2932
rect 39670 2887 39726 2896
rect 39488 2848 39540 2854
rect 39488 2790 39540 2796
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38384 2304 38436 2310
rect 38384 2246 38436 2252
rect 38396 1970 38424 2246
rect 38384 1964 38436 1970
rect 38384 1906 38436 1912
rect 38764 800 38792 2382
rect 39212 2304 39264 2310
rect 39212 2246 39264 2252
rect 39224 2106 39252 2246
rect 39212 2100 39264 2106
rect 39212 2042 39264 2048
rect 39500 800 39528 2790
rect 39868 2514 39896 2926
rect 40144 2774 40172 2994
rect 40236 2854 40264 3334
rect 40224 2848 40276 2854
rect 40224 2790 40276 2796
rect 40052 2746 40172 2774
rect 39856 2508 39908 2514
rect 39856 2450 39908 2456
rect 40052 2310 40080 2746
rect 40696 2446 40724 3402
rect 43352 3052 43404 3058
rect 43352 2994 43404 3000
rect 43168 2984 43220 2990
rect 43168 2926 43220 2932
rect 43180 2650 43208 2926
rect 43168 2644 43220 2650
rect 43168 2586 43220 2592
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 43272 2514 43300 2586
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 41144 2440 41196 2446
rect 41144 2382 41196 2388
rect 42708 2440 42760 2446
rect 43364 2428 43392 2994
rect 43628 2984 43680 2990
rect 43628 2926 43680 2932
rect 43640 2774 43668 2926
rect 43548 2746 43668 2774
rect 43444 2440 43496 2446
rect 43364 2400 43444 2428
rect 42708 2382 42760 2388
rect 43444 2382 43496 2388
rect 40040 2304 40092 2310
rect 40040 2246 40092 2252
rect 40408 2304 40460 2310
rect 40408 2246 40460 2252
rect 40420 1170 40448 2246
rect 40328 1142 40448 1170
rect 40328 800 40356 1142
rect 41156 800 41184 2382
rect 42720 800 42748 2382
rect 43548 800 43576 2746
rect 45480 2650 45508 3470
rect 46112 3460 46164 3466
rect 46112 3402 46164 3408
rect 46124 3346 46152 3402
rect 46388 3392 46440 3398
rect 46124 3318 46336 3346
rect 46388 3334 46440 3340
rect 46204 3188 46256 3194
rect 46204 3130 46256 3136
rect 46216 2854 46244 3130
rect 46308 2854 46336 3318
rect 46400 3058 46428 3334
rect 46388 3052 46440 3058
rect 46388 2994 46440 3000
rect 46204 2848 46256 2854
rect 46204 2790 46256 2796
rect 46296 2848 46348 2854
rect 46296 2790 46348 2796
rect 45468 2644 45520 2650
rect 45468 2586 45520 2592
rect 44088 2440 44140 2446
rect 44088 2382 44140 2388
rect 45100 2440 45152 2446
rect 45100 2382 45152 2388
rect 45928 2440 45980 2446
rect 45928 2382 45980 2388
rect 44100 2310 44128 2382
rect 44088 2304 44140 2310
rect 44088 2246 44140 2252
rect 44100 2106 44128 2246
rect 44088 2100 44140 2106
rect 44088 2042 44140 2048
rect 45112 800 45140 2382
rect 45940 800 45968 2382
rect 46492 1970 46520 3470
rect 47596 3074 47624 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 51908 3188 51960 3194
rect 51908 3130 51960 3136
rect 47596 3058 47808 3074
rect 47596 3052 47820 3058
rect 47596 3046 47768 3052
rect 47768 2994 47820 3000
rect 50620 3052 50672 3058
rect 50620 2994 50672 3000
rect 47584 2984 47636 2990
rect 47582 2952 47584 2961
rect 47636 2952 47638 2961
rect 47582 2887 47638 2896
rect 47780 2446 47808 2994
rect 50632 2961 50660 2994
rect 50618 2952 50674 2961
rect 50618 2887 50674 2896
rect 51920 2854 51948 3130
rect 52368 3052 52420 3058
rect 52368 2994 52420 3000
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 51908 2848 51960 2854
rect 51908 2790 51960 2796
rect 47492 2440 47544 2446
rect 47492 2382 47544 2388
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 49884 2440 49936 2446
rect 49884 2382 49936 2388
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 46860 2038 46888 2246
rect 46848 2032 46900 2038
rect 46848 1974 46900 1980
rect 46480 1964 46532 1970
rect 46480 1906 46532 1912
rect 47504 800 47532 2382
rect 47780 2106 47808 2382
rect 47768 2100 47820 2106
rect 47768 2042 47820 2048
rect 48332 800 48360 2382
rect 49896 800 49924 2382
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50724 800 50752 2790
rect 52276 2644 52328 2650
rect 52276 2586 52328 2592
rect 52288 2446 52316 2586
rect 52276 2440 52328 2446
rect 52276 2382 52328 2388
rect 52380 800 52408 2994
rect 52472 2650 52500 3470
rect 52840 3126 52868 3470
rect 53288 3460 53340 3466
rect 53288 3402 53340 3408
rect 53300 3194 53328 3402
rect 54956 3194 54984 37198
rect 55784 37126 55812 39200
rect 59268 37256 59320 37262
rect 59268 37198 59320 37204
rect 55772 37120 55824 37126
rect 55772 37062 55824 37068
rect 57336 18692 57388 18698
rect 57336 18634 57388 18640
rect 56968 3528 57020 3534
rect 56968 3470 57020 3476
rect 53288 3188 53340 3194
rect 53288 3130 53340 3136
rect 54944 3188 54996 3194
rect 54944 3130 54996 3136
rect 56980 3126 57008 3470
rect 52828 3120 52880 3126
rect 52828 3062 52880 3068
rect 56968 3120 57020 3126
rect 56968 3062 57020 3068
rect 53012 3052 53064 3058
rect 53012 2994 53064 3000
rect 56600 3052 56652 3058
rect 56784 3052 56836 3058
rect 56652 3012 56784 3040
rect 56600 2994 56652 3000
rect 56784 2994 56836 3000
rect 57152 3052 57204 3058
rect 57152 2994 57204 3000
rect 52460 2644 52512 2650
rect 52460 2586 52512 2592
rect 53024 2446 53052 2994
rect 54852 2984 54904 2990
rect 54852 2926 54904 2932
rect 53196 2644 53248 2650
rect 53196 2586 53248 2592
rect 53012 2440 53064 2446
rect 53012 2382 53064 2388
rect 53104 2440 53156 2446
rect 53104 2382 53156 2388
rect 53024 2310 53052 2382
rect 53012 2304 53064 2310
rect 53012 2246 53064 2252
rect 53116 800 53144 2382
rect 53208 2378 53236 2586
rect 54760 2440 54812 2446
rect 54760 2382 54812 2388
rect 53196 2372 53248 2378
rect 53196 2314 53248 2320
rect 54772 800 54800 2382
rect 54864 2038 54892 2926
rect 56612 2446 56640 2994
rect 55496 2440 55548 2446
rect 55496 2382 55548 2388
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 54852 2032 54904 2038
rect 54852 1974 54904 1980
rect 55508 800 55536 2382
rect 57164 800 57192 2994
rect 57348 2990 57376 18634
rect 57980 3936 58032 3942
rect 57980 3878 58032 3884
rect 57992 3194 58020 3878
rect 59280 3738 59308 37198
rect 59924 37126 59952 39200
rect 64064 37126 64092 39200
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 68204 37262 68232 39200
rect 76484 37330 76512 39200
rect 76472 37324 76524 37330
rect 76472 37266 76524 37272
rect 64144 37256 64196 37262
rect 64144 37198 64196 37204
rect 68192 37256 68244 37262
rect 68192 37198 68244 37204
rect 74632 37256 74684 37262
rect 74632 37198 74684 37204
rect 59912 37120 59964 37126
rect 59912 37062 59964 37068
rect 64052 37120 64104 37126
rect 64052 37062 64104 37068
rect 64156 36922 64184 37198
rect 64420 37120 64472 37126
rect 64420 37062 64472 37068
rect 64144 36916 64196 36922
rect 64144 36858 64196 36864
rect 64328 26784 64380 26790
rect 64328 26726 64380 26732
rect 64236 19780 64288 19786
rect 64236 19722 64288 19728
rect 64248 19514 64276 19722
rect 64236 19508 64288 19514
rect 64236 19450 64288 19456
rect 64052 5228 64104 5234
rect 64052 5170 64104 5176
rect 61660 5092 61712 5098
rect 61660 5034 61712 5040
rect 61672 4690 61700 5034
rect 63040 5024 63092 5030
rect 63040 4966 63092 4972
rect 61660 4684 61712 4690
rect 61660 4626 61712 4632
rect 63052 4622 63080 4966
rect 64064 4826 64092 5170
rect 63132 4820 63184 4826
rect 63132 4762 63184 4768
rect 64052 4820 64104 4826
rect 64052 4762 64104 4768
rect 63040 4616 63092 4622
rect 63040 4558 63092 4564
rect 63144 4078 63172 4762
rect 59452 4072 59504 4078
rect 59452 4014 59504 4020
rect 63132 4072 63184 4078
rect 63132 4014 63184 4020
rect 59268 3732 59320 3738
rect 59268 3674 59320 3680
rect 59464 3670 59492 4014
rect 62212 3936 62264 3942
rect 62212 3878 62264 3884
rect 59452 3664 59504 3670
rect 59452 3606 59504 3612
rect 62224 3534 62252 3878
rect 64340 3602 64368 26726
rect 64432 5370 64460 37062
rect 66352 36916 66404 36922
rect 66352 36858 66404 36864
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 66168 20460 66220 20466
rect 66168 20402 66220 20408
rect 64972 20324 65024 20330
rect 64972 20266 65024 20272
rect 64984 20058 65012 20266
rect 65432 20256 65484 20262
rect 65432 20198 65484 20204
rect 64972 20052 65024 20058
rect 64972 19994 65024 20000
rect 64880 19712 64932 19718
rect 64880 19654 64932 19660
rect 64892 19514 64920 19654
rect 64880 19508 64932 19514
rect 64880 19450 64932 19456
rect 65444 19378 65472 20198
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 65432 19372 65484 19378
rect 65432 19314 65484 19320
rect 66180 19310 66208 20402
rect 66168 19304 66220 19310
rect 66168 19246 66220 19252
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 64420 5364 64472 5370
rect 64420 5306 64472 5312
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 62212 3528 62264 3534
rect 62212 3470 62264 3476
rect 64052 3528 64104 3534
rect 64052 3470 64104 3476
rect 61752 3392 61804 3398
rect 61752 3334 61804 3340
rect 62396 3392 62448 3398
rect 62396 3334 62448 3340
rect 57980 3188 58032 3194
rect 57980 3130 58032 3136
rect 59544 3052 59596 3058
rect 59544 2994 59596 3000
rect 57336 2984 57388 2990
rect 57336 2926 57388 2932
rect 57440 2922 57652 2938
rect 57428 2916 57664 2922
rect 57480 2910 57612 2916
rect 57428 2858 57480 2864
rect 57612 2858 57664 2864
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 57900 800 57928 2382
rect 59556 800 59584 2994
rect 61764 2582 61792 3334
rect 62408 3194 62436 3334
rect 62396 3188 62448 3194
rect 62396 3130 62448 3136
rect 61844 3120 61896 3126
rect 61844 3062 61896 3068
rect 61752 2576 61804 2582
rect 61752 2518 61804 2524
rect 60372 2440 60424 2446
rect 60372 2382 60424 2388
rect 59820 2304 59872 2310
rect 59820 2246 59872 2252
rect 59832 2106 59860 2246
rect 59820 2100 59872 2106
rect 59820 2042 59872 2048
rect 60384 800 60412 2382
rect 61856 1578 61884 3062
rect 61936 3052 61988 3058
rect 61936 2994 61988 3000
rect 61948 2582 61976 2994
rect 62028 2848 62080 2854
rect 62028 2790 62080 2796
rect 62120 2848 62172 2854
rect 62120 2790 62172 2796
rect 62040 2582 62068 2790
rect 61936 2576 61988 2582
rect 61936 2518 61988 2524
rect 62028 2576 62080 2582
rect 62028 2518 62080 2524
rect 62132 2378 62160 2790
rect 64064 2582 64092 3470
rect 66364 3194 66392 36858
rect 68652 22568 68704 22574
rect 68652 22510 68704 22516
rect 68664 20602 68692 22510
rect 74644 20602 74672 37198
rect 84764 37126 84792 39200
rect 86868 37392 86920 37398
rect 86868 37334 86920 37340
rect 84844 37256 84896 37262
rect 84844 37198 84896 37204
rect 84752 37120 84804 37126
rect 84752 37062 84804 37068
rect 81014 37020 81322 37029
rect 81014 37018 81020 37020
rect 81076 37018 81100 37020
rect 81156 37018 81180 37020
rect 81236 37018 81260 37020
rect 81316 37018 81322 37020
rect 81076 36966 81078 37018
rect 81258 36966 81260 37018
rect 81014 36964 81020 36966
rect 81076 36964 81100 36966
rect 81156 36964 81180 36966
rect 81236 36964 81260 36966
rect 81316 36964 81322 36966
rect 81014 36955 81322 36964
rect 84856 36922 84884 37198
rect 84844 36916 84896 36922
rect 84844 36858 84896 36864
rect 86500 36100 86552 36106
rect 86500 36042 86552 36048
rect 81014 35932 81322 35941
rect 81014 35930 81020 35932
rect 81076 35930 81100 35932
rect 81156 35930 81180 35932
rect 81236 35930 81260 35932
rect 81316 35930 81322 35932
rect 81076 35878 81078 35930
rect 81258 35878 81260 35930
rect 81014 35876 81020 35878
rect 81076 35876 81100 35878
rect 81156 35876 81180 35878
rect 81236 35876 81260 35878
rect 81316 35876 81322 35878
rect 81014 35867 81322 35876
rect 81014 34844 81322 34853
rect 81014 34842 81020 34844
rect 81076 34842 81100 34844
rect 81156 34842 81180 34844
rect 81236 34842 81260 34844
rect 81316 34842 81322 34844
rect 81076 34790 81078 34842
rect 81258 34790 81260 34842
rect 81014 34788 81020 34790
rect 81076 34788 81100 34790
rect 81156 34788 81180 34790
rect 81236 34788 81260 34790
rect 81316 34788 81322 34790
rect 81014 34779 81322 34788
rect 81014 33756 81322 33765
rect 81014 33754 81020 33756
rect 81076 33754 81100 33756
rect 81156 33754 81180 33756
rect 81236 33754 81260 33756
rect 81316 33754 81322 33756
rect 81076 33702 81078 33754
rect 81258 33702 81260 33754
rect 81014 33700 81020 33702
rect 81076 33700 81100 33702
rect 81156 33700 81180 33702
rect 81236 33700 81260 33702
rect 81316 33700 81322 33702
rect 81014 33691 81322 33700
rect 81014 32668 81322 32677
rect 81014 32666 81020 32668
rect 81076 32666 81100 32668
rect 81156 32666 81180 32668
rect 81236 32666 81260 32668
rect 81316 32666 81322 32668
rect 81076 32614 81078 32666
rect 81258 32614 81260 32666
rect 81014 32612 81020 32614
rect 81076 32612 81100 32614
rect 81156 32612 81180 32614
rect 81236 32612 81260 32614
rect 81316 32612 81322 32614
rect 81014 32603 81322 32612
rect 81014 31580 81322 31589
rect 81014 31578 81020 31580
rect 81076 31578 81100 31580
rect 81156 31578 81180 31580
rect 81236 31578 81260 31580
rect 81316 31578 81322 31580
rect 81076 31526 81078 31578
rect 81258 31526 81260 31578
rect 81014 31524 81020 31526
rect 81076 31524 81100 31526
rect 81156 31524 81180 31526
rect 81236 31524 81260 31526
rect 81316 31524 81322 31526
rect 81014 31515 81322 31524
rect 81014 30492 81322 30501
rect 81014 30490 81020 30492
rect 81076 30490 81100 30492
rect 81156 30490 81180 30492
rect 81236 30490 81260 30492
rect 81316 30490 81322 30492
rect 81076 30438 81078 30490
rect 81258 30438 81260 30490
rect 81014 30436 81020 30438
rect 81076 30436 81100 30438
rect 81156 30436 81180 30438
rect 81236 30436 81260 30438
rect 81316 30436 81322 30438
rect 81014 30427 81322 30436
rect 81014 29404 81322 29413
rect 81014 29402 81020 29404
rect 81076 29402 81100 29404
rect 81156 29402 81180 29404
rect 81236 29402 81260 29404
rect 81316 29402 81322 29404
rect 81076 29350 81078 29402
rect 81258 29350 81260 29402
rect 81014 29348 81020 29350
rect 81076 29348 81100 29350
rect 81156 29348 81180 29350
rect 81236 29348 81260 29350
rect 81316 29348 81322 29350
rect 81014 29339 81322 29348
rect 81014 28316 81322 28325
rect 81014 28314 81020 28316
rect 81076 28314 81100 28316
rect 81156 28314 81180 28316
rect 81236 28314 81260 28316
rect 81316 28314 81322 28316
rect 81076 28262 81078 28314
rect 81258 28262 81260 28314
rect 81014 28260 81020 28262
rect 81076 28260 81100 28262
rect 81156 28260 81180 28262
rect 81236 28260 81260 28262
rect 81316 28260 81322 28262
rect 81014 28251 81322 28260
rect 81014 27228 81322 27237
rect 81014 27226 81020 27228
rect 81076 27226 81100 27228
rect 81156 27226 81180 27228
rect 81236 27226 81260 27228
rect 81316 27226 81322 27228
rect 81076 27174 81078 27226
rect 81258 27174 81260 27226
rect 81014 27172 81020 27174
rect 81076 27172 81100 27174
rect 81156 27172 81180 27174
rect 81236 27172 81260 27174
rect 81316 27172 81322 27174
rect 81014 27163 81322 27172
rect 81014 26140 81322 26149
rect 81014 26138 81020 26140
rect 81076 26138 81100 26140
rect 81156 26138 81180 26140
rect 81236 26138 81260 26140
rect 81316 26138 81322 26140
rect 81076 26086 81078 26138
rect 81258 26086 81260 26138
rect 81014 26084 81020 26086
rect 81076 26084 81100 26086
rect 81156 26084 81180 26086
rect 81236 26084 81260 26086
rect 81316 26084 81322 26086
rect 81014 26075 81322 26084
rect 81014 25052 81322 25061
rect 81014 25050 81020 25052
rect 81076 25050 81100 25052
rect 81156 25050 81180 25052
rect 81236 25050 81260 25052
rect 81316 25050 81322 25052
rect 81076 24998 81078 25050
rect 81258 24998 81260 25050
rect 81014 24996 81020 24998
rect 81076 24996 81100 24998
rect 81156 24996 81180 24998
rect 81236 24996 81260 24998
rect 81316 24996 81322 24998
rect 81014 24987 81322 24996
rect 81014 23964 81322 23973
rect 81014 23962 81020 23964
rect 81076 23962 81100 23964
rect 81156 23962 81180 23964
rect 81236 23962 81260 23964
rect 81316 23962 81322 23964
rect 81076 23910 81078 23962
rect 81258 23910 81260 23962
rect 81014 23908 81020 23910
rect 81076 23908 81100 23910
rect 81156 23908 81180 23910
rect 81236 23908 81260 23910
rect 81316 23908 81322 23910
rect 81014 23899 81322 23908
rect 81014 22876 81322 22885
rect 81014 22874 81020 22876
rect 81076 22874 81100 22876
rect 81156 22874 81180 22876
rect 81236 22874 81260 22876
rect 81316 22874 81322 22876
rect 81076 22822 81078 22874
rect 81258 22822 81260 22874
rect 81014 22820 81020 22822
rect 81076 22820 81100 22822
rect 81156 22820 81180 22822
rect 81236 22820 81260 22822
rect 81316 22820 81322 22822
rect 81014 22811 81322 22820
rect 81014 21788 81322 21797
rect 81014 21786 81020 21788
rect 81076 21786 81100 21788
rect 81156 21786 81180 21788
rect 81236 21786 81260 21788
rect 81316 21786 81322 21788
rect 81076 21734 81078 21786
rect 81258 21734 81260 21786
rect 81014 21732 81020 21734
rect 81076 21732 81100 21734
rect 81156 21732 81180 21734
rect 81236 21732 81260 21734
rect 81316 21732 81322 21734
rect 81014 21723 81322 21732
rect 77116 20800 77168 20806
rect 77116 20742 77168 20748
rect 68652 20596 68704 20602
rect 68652 20538 68704 20544
rect 69296 20596 69348 20602
rect 69296 20538 69348 20544
rect 70400 20596 70452 20602
rect 70400 20538 70452 20544
rect 74632 20596 74684 20602
rect 74632 20538 74684 20544
rect 68836 20460 68888 20466
rect 68836 20402 68888 20408
rect 68848 20058 68876 20402
rect 69308 20398 69336 20538
rect 70412 20398 70440 20538
rect 70676 20528 70728 20534
rect 70676 20470 70728 20476
rect 69296 20392 69348 20398
rect 69296 20334 69348 20340
rect 69388 20392 69440 20398
rect 69388 20334 69440 20340
rect 70400 20392 70452 20398
rect 70400 20334 70452 20340
rect 69020 20256 69072 20262
rect 69020 20198 69072 20204
rect 68836 20052 68888 20058
rect 68836 19994 68888 20000
rect 68376 19916 68428 19922
rect 68376 19858 68428 19864
rect 68388 19310 68416 19858
rect 69032 19854 69060 20198
rect 69400 19922 69428 20334
rect 70032 20256 70084 20262
rect 70032 20198 70084 20204
rect 69388 19916 69440 19922
rect 69388 19858 69440 19864
rect 69020 19848 69072 19854
rect 69020 19790 69072 19796
rect 68376 19304 68428 19310
rect 68376 19246 68428 19252
rect 68560 5024 68612 5030
rect 68560 4966 68612 4972
rect 68572 4622 68600 4966
rect 69204 4820 69256 4826
rect 69204 4762 69256 4768
rect 68560 4616 68612 4622
rect 68560 4558 68612 4564
rect 69216 4078 69244 4762
rect 69400 4554 69428 19858
rect 70044 19378 70072 20198
rect 70032 19372 70084 19378
rect 70032 19314 70084 19320
rect 70688 19174 70716 20470
rect 74908 20460 74960 20466
rect 74908 20402 74960 20408
rect 74724 20392 74776 20398
rect 74724 20334 74776 20340
rect 73620 20256 73672 20262
rect 73620 20198 73672 20204
rect 73632 19854 73660 20198
rect 73620 19848 73672 19854
rect 73620 19790 73672 19796
rect 70860 19712 70912 19718
rect 70860 19654 70912 19660
rect 70872 19378 70900 19654
rect 73896 19508 73948 19514
rect 73896 19450 73948 19456
rect 70860 19372 70912 19378
rect 70860 19314 70912 19320
rect 70676 19168 70728 19174
rect 70676 19110 70728 19116
rect 73908 16574 73936 19450
rect 73908 16546 74028 16574
rect 70492 15360 70544 15366
rect 70492 15302 70544 15308
rect 70504 5370 70532 15302
rect 70492 5364 70544 5370
rect 70492 5306 70544 5312
rect 70124 5228 70176 5234
rect 70124 5170 70176 5176
rect 70136 4826 70164 5170
rect 73436 5024 73488 5030
rect 73436 4966 73488 4972
rect 70124 4820 70176 4826
rect 70124 4762 70176 4768
rect 73448 4622 73476 4966
rect 74000 4690 74028 16546
rect 74448 5296 74500 5302
rect 74448 5238 74500 5244
rect 73988 4684 74040 4690
rect 73988 4626 74040 4632
rect 73436 4616 73488 4622
rect 73436 4558 73488 4564
rect 69388 4548 69440 4554
rect 69388 4490 69440 4496
rect 74460 4486 74488 5238
rect 73896 4480 73948 4486
rect 73896 4422 73948 4428
rect 74448 4480 74500 4486
rect 74448 4422 74500 4428
rect 73908 4146 73936 4422
rect 73896 4140 73948 4146
rect 73896 4082 73948 4088
rect 73988 4140 74040 4146
rect 73988 4082 74040 4088
rect 69204 4072 69256 4078
rect 69204 4014 69256 4020
rect 68376 4004 68428 4010
rect 68376 3946 68428 3952
rect 68192 3936 68244 3942
rect 68192 3878 68244 3884
rect 66812 3528 66864 3534
rect 66812 3470 66864 3476
rect 66352 3188 66404 3194
rect 66352 3130 66404 3136
rect 66260 3052 66312 3058
rect 66260 2994 66312 3000
rect 65156 2848 65208 2854
rect 65156 2790 65208 2796
rect 64052 2576 64104 2582
rect 64052 2518 64104 2524
rect 62672 2508 62724 2514
rect 62672 2450 62724 2456
rect 62684 2417 62712 2450
rect 64328 2440 64380 2446
rect 62670 2408 62726 2417
rect 62120 2372 62172 2378
rect 64328 2382 64380 2388
rect 62670 2343 62726 2352
rect 62764 2372 62816 2378
rect 62120 2314 62172 2320
rect 62764 2314 62816 2320
rect 61856 1550 61976 1578
rect 61948 800 61976 1550
rect 62776 800 62804 2314
rect 64340 800 64368 2382
rect 65168 800 65196 2790
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66272 2582 66300 2994
rect 65800 2576 65852 2582
rect 65800 2518 65852 2524
rect 66260 2576 66312 2582
rect 66260 2518 66312 2524
rect 65812 2446 65840 2518
rect 66824 2514 66852 3470
rect 68204 3058 68232 3878
rect 68388 3194 68416 3946
rect 73620 3936 73672 3942
rect 73620 3878 73672 3884
rect 68836 3528 68888 3534
rect 68836 3470 68888 3476
rect 68376 3188 68428 3194
rect 68376 3130 68428 3136
rect 68192 3052 68244 3058
rect 68192 2994 68244 3000
rect 68652 2984 68704 2990
rect 68652 2926 68704 2932
rect 67548 2576 67600 2582
rect 67548 2518 67600 2524
rect 66812 2508 66864 2514
rect 66812 2450 66864 2456
rect 65800 2440 65852 2446
rect 65706 2408 65762 2417
rect 65800 2382 65852 2388
rect 66720 2440 66772 2446
rect 66720 2382 66772 2388
rect 65706 2343 65762 2352
rect 65720 2310 65748 2343
rect 65708 2304 65760 2310
rect 65708 2246 65760 2252
rect 66732 800 66760 2382
rect 67560 800 67588 2518
rect 68664 2446 68692 2926
rect 68848 2514 68876 3470
rect 73632 3058 73660 3878
rect 74000 3670 74028 4082
rect 74736 4078 74764 20334
rect 74920 20058 74948 20402
rect 74908 20052 74960 20058
rect 74908 19994 74960 20000
rect 77128 6458 77156 20742
rect 81014 20700 81322 20709
rect 81014 20698 81020 20700
rect 81076 20698 81100 20700
rect 81156 20698 81180 20700
rect 81236 20698 81260 20700
rect 81316 20698 81322 20700
rect 81076 20646 81078 20698
rect 81258 20646 81260 20698
rect 81014 20644 81020 20646
rect 81076 20644 81100 20646
rect 81156 20644 81180 20646
rect 81236 20644 81260 20646
rect 81316 20644 81322 20646
rect 81014 20635 81322 20644
rect 81014 19612 81322 19621
rect 81014 19610 81020 19612
rect 81076 19610 81100 19612
rect 81156 19610 81180 19612
rect 81236 19610 81260 19612
rect 81316 19610 81322 19612
rect 81076 19558 81078 19610
rect 81258 19558 81260 19610
rect 81014 19556 81020 19558
rect 81076 19556 81100 19558
rect 81156 19556 81180 19558
rect 81236 19556 81260 19558
rect 81316 19556 81322 19558
rect 81014 19547 81322 19556
rect 81014 18524 81322 18533
rect 81014 18522 81020 18524
rect 81076 18522 81100 18524
rect 81156 18522 81180 18524
rect 81236 18522 81260 18524
rect 81316 18522 81322 18524
rect 81076 18470 81078 18522
rect 81258 18470 81260 18522
rect 81014 18468 81020 18470
rect 81076 18468 81100 18470
rect 81156 18468 81180 18470
rect 81236 18468 81260 18470
rect 81316 18468 81322 18470
rect 81014 18459 81322 18468
rect 81014 17436 81322 17445
rect 81014 17434 81020 17436
rect 81076 17434 81100 17436
rect 81156 17434 81180 17436
rect 81236 17434 81260 17436
rect 81316 17434 81322 17436
rect 81076 17382 81078 17434
rect 81258 17382 81260 17434
rect 81014 17380 81020 17382
rect 81076 17380 81100 17382
rect 81156 17380 81180 17382
rect 81236 17380 81260 17382
rect 81316 17380 81322 17382
rect 81014 17371 81322 17380
rect 81014 16348 81322 16357
rect 81014 16346 81020 16348
rect 81076 16346 81100 16348
rect 81156 16346 81180 16348
rect 81236 16346 81260 16348
rect 81316 16346 81322 16348
rect 81076 16294 81078 16346
rect 81258 16294 81260 16346
rect 81014 16292 81020 16294
rect 81076 16292 81100 16294
rect 81156 16292 81180 16294
rect 81236 16292 81260 16294
rect 81316 16292 81322 16294
rect 81014 16283 81322 16292
rect 81014 15260 81322 15269
rect 81014 15258 81020 15260
rect 81076 15258 81100 15260
rect 81156 15258 81180 15260
rect 81236 15258 81260 15260
rect 81316 15258 81322 15260
rect 81076 15206 81078 15258
rect 81258 15206 81260 15258
rect 81014 15204 81020 15206
rect 81076 15204 81100 15206
rect 81156 15204 81180 15206
rect 81236 15204 81260 15206
rect 81316 15204 81322 15206
rect 81014 15195 81322 15204
rect 81014 14172 81322 14181
rect 81014 14170 81020 14172
rect 81076 14170 81100 14172
rect 81156 14170 81180 14172
rect 81236 14170 81260 14172
rect 81316 14170 81322 14172
rect 81076 14118 81078 14170
rect 81258 14118 81260 14170
rect 81014 14116 81020 14118
rect 81076 14116 81100 14118
rect 81156 14116 81180 14118
rect 81236 14116 81260 14118
rect 81316 14116 81322 14118
rect 81014 14107 81322 14116
rect 81014 13084 81322 13093
rect 81014 13082 81020 13084
rect 81076 13082 81100 13084
rect 81156 13082 81180 13084
rect 81236 13082 81260 13084
rect 81316 13082 81322 13084
rect 81076 13030 81078 13082
rect 81258 13030 81260 13082
rect 81014 13028 81020 13030
rect 81076 13028 81100 13030
rect 81156 13028 81180 13030
rect 81236 13028 81260 13030
rect 81316 13028 81322 13030
rect 81014 13019 81322 13028
rect 81014 11996 81322 12005
rect 81014 11994 81020 11996
rect 81076 11994 81100 11996
rect 81156 11994 81180 11996
rect 81236 11994 81260 11996
rect 81316 11994 81322 11996
rect 81076 11942 81078 11994
rect 81258 11942 81260 11994
rect 81014 11940 81020 11942
rect 81076 11940 81100 11942
rect 81156 11940 81180 11942
rect 81236 11940 81260 11942
rect 81316 11940 81322 11942
rect 81014 11931 81322 11940
rect 81014 10908 81322 10917
rect 81014 10906 81020 10908
rect 81076 10906 81100 10908
rect 81156 10906 81180 10908
rect 81236 10906 81260 10908
rect 81316 10906 81322 10908
rect 81076 10854 81078 10906
rect 81258 10854 81260 10906
rect 81014 10852 81020 10854
rect 81076 10852 81100 10854
rect 81156 10852 81180 10854
rect 81236 10852 81260 10854
rect 81316 10852 81322 10854
rect 81014 10843 81322 10852
rect 81014 9820 81322 9829
rect 81014 9818 81020 9820
rect 81076 9818 81100 9820
rect 81156 9818 81180 9820
rect 81236 9818 81260 9820
rect 81316 9818 81322 9820
rect 81076 9766 81078 9818
rect 81258 9766 81260 9818
rect 81014 9764 81020 9766
rect 81076 9764 81100 9766
rect 81156 9764 81180 9766
rect 81236 9764 81260 9766
rect 81316 9764 81322 9766
rect 81014 9755 81322 9764
rect 81014 8732 81322 8741
rect 81014 8730 81020 8732
rect 81076 8730 81100 8732
rect 81156 8730 81180 8732
rect 81236 8730 81260 8732
rect 81316 8730 81322 8732
rect 81076 8678 81078 8730
rect 81258 8678 81260 8730
rect 81014 8676 81020 8678
rect 81076 8676 81100 8678
rect 81156 8676 81180 8678
rect 81236 8676 81260 8678
rect 81316 8676 81322 8678
rect 81014 8667 81322 8676
rect 81014 7644 81322 7653
rect 81014 7642 81020 7644
rect 81076 7642 81100 7644
rect 81156 7642 81180 7644
rect 81236 7642 81260 7644
rect 81316 7642 81322 7644
rect 81076 7590 81078 7642
rect 81258 7590 81260 7642
rect 81014 7588 81020 7590
rect 81076 7588 81100 7590
rect 81156 7588 81180 7590
rect 81236 7588 81260 7590
rect 81316 7588 81322 7590
rect 81014 7579 81322 7588
rect 81014 6556 81322 6565
rect 81014 6554 81020 6556
rect 81076 6554 81100 6556
rect 81156 6554 81180 6556
rect 81236 6554 81260 6556
rect 81316 6554 81322 6556
rect 81076 6502 81078 6554
rect 81258 6502 81260 6554
rect 81014 6500 81020 6502
rect 81076 6500 81100 6502
rect 81156 6500 81180 6502
rect 81236 6500 81260 6502
rect 81316 6500 81322 6502
rect 81014 6491 81322 6500
rect 77116 6452 77168 6458
rect 77116 6394 77168 6400
rect 76932 6316 76984 6322
rect 76932 6258 76984 6264
rect 76012 6112 76064 6118
rect 76012 6054 76064 6060
rect 76024 5710 76052 6054
rect 75920 5704 75972 5710
rect 75920 5646 75972 5652
rect 76012 5704 76064 5710
rect 76012 5646 76064 5652
rect 75932 4758 75960 5646
rect 76944 5574 76972 6258
rect 77208 6248 77260 6254
rect 77208 6190 77260 6196
rect 76932 5568 76984 5574
rect 76932 5510 76984 5516
rect 76944 4826 76972 5510
rect 77220 5166 77248 6190
rect 81014 5468 81322 5477
rect 81014 5466 81020 5468
rect 81076 5466 81100 5468
rect 81156 5466 81180 5468
rect 81236 5466 81260 5468
rect 81316 5466 81322 5468
rect 81076 5414 81078 5466
rect 81258 5414 81260 5466
rect 81014 5412 81020 5414
rect 81076 5412 81100 5414
rect 81156 5412 81180 5414
rect 81236 5412 81260 5414
rect 81316 5412 81322 5414
rect 81014 5403 81322 5412
rect 77208 5160 77260 5166
rect 77208 5102 77260 5108
rect 77300 5092 77352 5098
rect 77300 5034 77352 5040
rect 76932 4820 76984 4826
rect 76932 4762 76984 4768
rect 75920 4752 75972 4758
rect 75920 4694 75972 4700
rect 75932 4554 75960 4694
rect 75920 4548 75972 4554
rect 75920 4490 75972 4496
rect 76748 4548 76800 4554
rect 76748 4490 76800 4496
rect 74724 4072 74776 4078
rect 74724 4014 74776 4020
rect 73988 3664 74040 3670
rect 73988 3606 74040 3612
rect 73896 3528 73948 3534
rect 73896 3470 73948 3476
rect 73620 3052 73672 3058
rect 73620 2994 73672 3000
rect 73712 3052 73764 3058
rect 73712 2994 73764 3000
rect 70768 2984 70820 2990
rect 70768 2926 70820 2932
rect 68836 2508 68888 2514
rect 70032 2508 70084 2514
rect 68836 2450 68888 2456
rect 69952 2468 70032 2496
rect 68652 2440 68704 2446
rect 68652 2382 68704 2388
rect 69112 1420 69164 1426
rect 69112 1362 69164 1368
rect 69124 800 69152 1362
rect 69952 800 69980 2468
rect 70032 2450 70084 2456
rect 70124 2440 70176 2446
rect 70124 2382 70176 2388
rect 70136 1426 70164 2382
rect 70780 2378 70808 2926
rect 73724 2582 73752 2994
rect 73712 2576 73764 2582
rect 73712 2518 73764 2524
rect 71504 2440 71556 2446
rect 71504 2382 71556 2388
rect 72332 2440 72384 2446
rect 72332 2382 72384 2388
rect 70768 2372 70820 2378
rect 70768 2314 70820 2320
rect 70124 1420 70176 1426
rect 70124 1362 70176 1368
rect 71516 800 71544 2382
rect 72344 800 72372 2382
rect 73908 800 73936 3470
rect 74000 2922 74028 3606
rect 74540 3392 74592 3398
rect 74540 3334 74592 3340
rect 73988 2916 74040 2922
rect 73988 2858 74040 2864
rect 74552 2514 74580 3334
rect 76760 3058 76788 4490
rect 77312 4282 77340 5034
rect 86224 4752 86276 4758
rect 86224 4694 86276 4700
rect 78588 4480 78640 4486
rect 78588 4422 78640 4428
rect 77300 4276 77352 4282
rect 77300 4218 77352 4224
rect 77312 4146 77340 4218
rect 77300 4140 77352 4146
rect 77300 4082 77352 4088
rect 78600 3602 78628 4422
rect 81014 4380 81322 4389
rect 81014 4378 81020 4380
rect 81076 4378 81100 4380
rect 81156 4378 81180 4380
rect 81236 4378 81260 4380
rect 81316 4378 81322 4380
rect 81076 4326 81078 4378
rect 81258 4326 81260 4378
rect 81014 4324 81020 4326
rect 81076 4324 81100 4326
rect 81156 4324 81180 4326
rect 81236 4324 81260 4326
rect 81316 4324 81322 4326
rect 81014 4315 81322 4324
rect 79140 3732 79192 3738
rect 79140 3674 79192 3680
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 79152 3126 79180 3674
rect 86236 3602 86264 4694
rect 86316 4276 86368 4282
rect 86316 4218 86368 4224
rect 86328 4146 86356 4218
rect 86316 4140 86368 4146
rect 86316 4082 86368 4088
rect 86512 4078 86540 36042
rect 86500 4072 86552 4078
rect 86500 4014 86552 4020
rect 86512 3942 86540 4014
rect 86316 3936 86368 3942
rect 86316 3878 86368 3884
rect 86500 3936 86552 3942
rect 86500 3878 86552 3884
rect 86224 3596 86276 3602
rect 86224 3538 86276 3544
rect 86328 3534 86356 3878
rect 83556 3528 83608 3534
rect 83556 3470 83608 3476
rect 86316 3528 86368 3534
rect 86316 3470 86368 3476
rect 81014 3292 81322 3301
rect 81014 3290 81020 3292
rect 81076 3290 81100 3292
rect 81156 3290 81180 3292
rect 81236 3290 81260 3292
rect 81316 3290 81322 3292
rect 81076 3238 81078 3290
rect 81258 3238 81260 3290
rect 81014 3236 81020 3238
rect 81076 3236 81100 3238
rect 81156 3236 81180 3238
rect 81236 3236 81260 3238
rect 81316 3236 81322 3238
rect 81014 3227 81322 3236
rect 83568 3194 83596 3470
rect 83648 3392 83700 3398
rect 83648 3334 83700 3340
rect 83556 3188 83608 3194
rect 83556 3130 83608 3136
rect 79140 3120 79192 3126
rect 79140 3062 79192 3068
rect 83660 3058 83688 3334
rect 86880 3058 86908 37334
rect 92020 37324 92072 37330
rect 92020 37266 92072 37272
rect 88708 36576 88760 36582
rect 88708 36518 88760 36524
rect 87604 4140 87656 4146
rect 87604 4082 87656 4088
rect 87236 4004 87288 4010
rect 87236 3946 87288 3952
rect 87248 3738 87276 3946
rect 87236 3732 87288 3738
rect 87236 3674 87288 3680
rect 87616 3602 87644 4082
rect 87604 3596 87656 3602
rect 87604 3538 87656 3544
rect 88720 3534 88748 36518
rect 90272 35080 90324 35086
rect 90272 35022 90324 35028
rect 89076 3936 89128 3942
rect 89076 3878 89128 3884
rect 88708 3528 88760 3534
rect 88708 3470 88760 3476
rect 87696 3460 87748 3466
rect 87696 3402 87748 3408
rect 76288 3052 76340 3058
rect 76288 2994 76340 3000
rect 76748 3052 76800 3058
rect 76748 2994 76800 3000
rect 83648 3052 83700 3058
rect 83648 2994 83700 3000
rect 85948 3052 86000 3058
rect 85948 2994 86000 3000
rect 86868 3052 86920 3058
rect 86868 2994 86920 3000
rect 74632 2848 74684 2854
rect 74632 2790 74684 2796
rect 74724 2848 74776 2854
rect 74724 2790 74776 2796
rect 74540 2508 74592 2514
rect 74540 2450 74592 2456
rect 74644 1494 74672 2790
rect 74632 1488 74684 1494
rect 74632 1430 74684 1436
rect 74736 800 74764 2790
rect 76104 2304 76156 2310
rect 76104 2246 76156 2252
rect 76116 2038 76144 2246
rect 76104 2032 76156 2038
rect 76104 1974 76156 1980
rect 76300 800 76328 2994
rect 79968 2984 80020 2990
rect 79968 2926 80020 2932
rect 76380 2848 76432 2854
rect 76380 2790 76432 2796
rect 77116 2848 77168 2854
rect 77116 2790 77168 2796
rect 76392 2514 76420 2790
rect 76380 2508 76432 2514
rect 76380 2450 76432 2456
rect 77128 800 77156 2790
rect 79980 2582 80008 2926
rect 81900 2848 81952 2854
rect 81900 2790 81952 2796
rect 79048 2576 79100 2582
rect 79048 2518 79100 2524
rect 79968 2576 80020 2582
rect 79968 2518 80020 2524
rect 78680 2440 78732 2446
rect 78680 2382 78732 2388
rect 78692 800 78720 2382
rect 79060 2378 79088 2518
rect 79508 2440 79560 2446
rect 79508 2382 79560 2388
rect 81348 2440 81400 2446
rect 81348 2382 81400 2388
rect 79048 2372 79100 2378
rect 79048 2314 79100 2320
rect 79140 2304 79192 2310
rect 79140 2246 79192 2252
rect 79152 1630 79180 2246
rect 79140 1624 79192 1630
rect 79140 1566 79192 1572
rect 79520 800 79548 2382
rect 81014 2204 81322 2213
rect 81014 2202 81020 2204
rect 81076 2202 81100 2204
rect 81156 2202 81180 2204
rect 81236 2202 81260 2204
rect 81316 2202 81322 2204
rect 81076 2150 81078 2202
rect 81258 2150 81260 2202
rect 81014 2148 81020 2150
rect 81076 2148 81100 2150
rect 81156 2148 81180 2150
rect 81236 2148 81260 2150
rect 81316 2148 81322 2150
rect 81014 2139 81322 2148
rect 81360 1306 81388 2382
rect 81176 1278 81388 1306
rect 81176 800 81204 1278
rect 81912 800 81940 2790
rect 85396 2644 85448 2650
rect 85396 2586 85448 2592
rect 81992 2508 82044 2514
rect 81992 2450 82044 2456
rect 84844 2508 84896 2514
rect 84844 2450 84896 2456
rect 82004 1970 82032 2450
rect 83556 2440 83608 2446
rect 83556 2382 83608 2388
rect 84292 2440 84344 2446
rect 84292 2382 84344 2388
rect 81992 1964 82044 1970
rect 81992 1906 82044 1912
rect 83568 800 83596 2382
rect 84304 800 84332 2382
rect 84856 1970 84884 2450
rect 84844 1964 84896 1970
rect 84844 1906 84896 1912
rect 85408 1902 85436 2586
rect 85396 1896 85448 1902
rect 85396 1838 85448 1844
rect 85960 800 85988 2994
rect 87708 2854 87736 3402
rect 88156 3052 88208 3058
rect 88156 2994 88208 3000
rect 87696 2848 87748 2854
rect 87696 2790 87748 2796
rect 87972 2848 88024 2854
rect 87972 2790 88024 2796
rect 87984 2446 88012 2790
rect 88168 2650 88196 2994
rect 88156 2644 88208 2650
rect 88156 2586 88208 2592
rect 87972 2440 88024 2446
rect 87972 2382 88024 2388
rect 88156 2440 88208 2446
rect 88156 2382 88208 2388
rect 86776 2304 86828 2310
rect 86776 2246 86828 2252
rect 86788 1970 86816 2246
rect 86776 1964 86828 1970
rect 86776 1906 86828 1912
rect 88168 1426 88196 2382
rect 86684 1420 86736 1426
rect 86684 1362 86736 1368
rect 88156 1420 88208 1426
rect 88156 1362 88208 1368
rect 88340 1420 88392 1426
rect 88340 1362 88392 1368
rect 86696 800 86724 1362
rect 88352 800 88380 1362
rect 89088 800 89116 3878
rect 89628 3392 89680 3398
rect 89628 3334 89680 3340
rect 89640 3126 89668 3334
rect 89628 3120 89680 3126
rect 89628 3062 89680 3068
rect 89352 3052 89404 3058
rect 89352 2994 89404 3000
rect 89364 2854 89392 2994
rect 90284 2854 90312 35022
rect 92032 5370 92060 37266
rect 93044 37262 93072 39200
rect 96374 37564 96682 37573
rect 96374 37562 96380 37564
rect 96436 37562 96460 37564
rect 96516 37562 96540 37564
rect 96596 37562 96620 37564
rect 96676 37562 96682 37564
rect 96436 37510 96438 37562
rect 96618 37510 96620 37562
rect 96374 37508 96380 37510
rect 96436 37508 96460 37510
rect 96516 37508 96540 37510
rect 96596 37508 96620 37510
rect 96676 37508 96682 37510
rect 96374 37499 96682 37508
rect 93032 37256 93084 37262
rect 93032 37198 93084 37204
rect 109604 37126 109632 39200
rect 117226 39199 117282 39208
rect 117870 39200 117926 40000
rect 109684 37256 109736 37262
rect 109684 37198 109736 37204
rect 109592 37120 109644 37126
rect 109592 37062 109644 37068
rect 101772 36848 101824 36854
rect 101772 36790 101824 36796
rect 92112 36780 92164 36786
rect 92112 36722 92164 36728
rect 92020 5364 92072 5370
rect 92020 5306 92072 5312
rect 91928 5228 91980 5234
rect 91928 5170 91980 5176
rect 91100 5024 91152 5030
rect 91100 4966 91152 4972
rect 90364 4548 90416 4554
rect 90364 4490 90416 4496
rect 90376 4282 90404 4490
rect 90364 4276 90416 4282
rect 90364 4218 90416 4224
rect 91112 4146 91140 4966
rect 91940 4826 91968 5170
rect 91928 4820 91980 4826
rect 91928 4762 91980 4768
rect 91100 4140 91152 4146
rect 91100 4082 91152 4088
rect 90732 4072 90784 4078
rect 90732 4014 90784 4020
rect 90548 3936 90600 3942
rect 90548 3878 90600 3884
rect 89352 2848 89404 2854
rect 89352 2790 89404 2796
rect 90272 2848 90324 2854
rect 90272 2790 90324 2796
rect 89444 2644 89496 2650
rect 89444 2586 89496 2592
rect 89456 2378 89484 2586
rect 90456 2508 90508 2514
rect 90456 2450 90508 2456
rect 89628 2440 89680 2446
rect 89628 2382 89680 2388
rect 89444 2372 89496 2378
rect 89444 2314 89496 2320
rect 89640 1426 89668 2382
rect 90468 1834 90496 2450
rect 90560 2446 90588 3878
rect 90640 2916 90692 2922
rect 90640 2858 90692 2864
rect 90652 2446 90680 2858
rect 90548 2440 90600 2446
rect 90548 2382 90600 2388
rect 90640 2440 90692 2446
rect 90640 2382 90692 2388
rect 90456 1828 90508 1834
rect 90456 1770 90508 1776
rect 89628 1420 89680 1426
rect 89628 1362 89680 1368
rect 90744 800 90772 4014
rect 91652 4004 91704 4010
rect 91652 3946 91704 3952
rect 91664 3754 91692 3946
rect 91572 3738 91692 3754
rect 91560 3732 91692 3738
rect 91612 3726 91692 3732
rect 91744 3732 91796 3738
rect 91560 3674 91612 3680
rect 91744 3674 91796 3680
rect 91756 3602 91784 3674
rect 91940 3602 91968 4762
rect 91744 3596 91796 3602
rect 91744 3538 91796 3544
rect 91928 3596 91980 3602
rect 91928 3538 91980 3544
rect 91652 3528 91704 3534
rect 91652 3470 91704 3476
rect 91192 3392 91244 3398
rect 91192 3334 91244 3340
rect 91204 3058 91232 3334
rect 91192 3052 91244 3058
rect 91192 2994 91244 3000
rect 91664 2514 91692 3470
rect 91744 3460 91796 3466
rect 91744 3402 91796 3408
rect 91836 3460 91888 3466
rect 91836 3402 91888 3408
rect 91756 2922 91784 3402
rect 91744 2916 91796 2922
rect 91744 2858 91796 2864
rect 91848 2650 91876 3402
rect 92020 3052 92072 3058
rect 92020 2994 92072 3000
rect 91836 2644 91888 2650
rect 91836 2586 91888 2592
rect 91928 2644 91980 2650
rect 91928 2586 91980 2592
rect 91652 2508 91704 2514
rect 91652 2450 91704 2456
rect 91572 870 91692 898
rect 91572 800 91600 870
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4342 0 4398 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8298 0 8354 800
rect 9126 0 9182 800
rect 9954 0 10010 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12346 0 12402 800
rect 13174 0 13230 800
rect 13910 0 13966 800
rect 14738 0 14794 800
rect 15566 0 15622 800
rect 16302 0 16358 800
rect 17130 0 17186 800
rect 17958 0 18014 800
rect 18694 0 18750 800
rect 19522 0 19578 800
rect 20350 0 20406 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22742 0 22798 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25134 0 25190 800
rect 25962 0 26018 800
rect 26698 0 26754 800
rect 27526 0 27582 800
rect 28354 0 28410 800
rect 29090 0 29146 800
rect 29918 0 29974 800
rect 30746 0 30802 800
rect 31574 0 31630 800
rect 32310 0 32366 800
rect 33138 0 33194 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35530 0 35586 800
rect 36358 0 36414 800
rect 37094 0 37150 800
rect 37922 0 37978 800
rect 38750 0 38806 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45098 0 45154 800
rect 45926 0 45982 800
rect 46754 0 46810 800
rect 47490 0 47546 800
rect 48318 0 48374 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50710 0 50766 800
rect 51538 0 51594 800
rect 52366 0 52422 800
rect 53102 0 53158 800
rect 53930 0 53986 800
rect 54758 0 54814 800
rect 55494 0 55550 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 57886 0 57942 800
rect 58714 0 58770 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61106 0 61162 800
rect 61934 0 61990 800
rect 62762 0 62818 800
rect 63498 0 63554 800
rect 64326 0 64382 800
rect 65154 0 65210 800
rect 65890 0 65946 800
rect 66718 0 66774 800
rect 67546 0 67602 800
rect 68282 0 68338 800
rect 69110 0 69166 800
rect 69938 0 69994 800
rect 70766 0 70822 800
rect 71502 0 71558 800
rect 72330 0 72386 800
rect 73158 0 73214 800
rect 73894 0 73950 800
rect 74722 0 74778 800
rect 75550 0 75606 800
rect 76286 0 76342 800
rect 77114 0 77170 800
rect 77942 0 77998 800
rect 78678 0 78734 800
rect 79506 0 79562 800
rect 80334 0 80390 800
rect 81162 0 81218 800
rect 81898 0 81954 800
rect 82726 0 82782 800
rect 83554 0 83610 800
rect 84290 0 84346 800
rect 85118 0 85174 800
rect 85946 0 86002 800
rect 86682 0 86738 800
rect 87510 0 87566 800
rect 88338 0 88394 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 91664 762 91692 870
rect 91940 762 91968 2586
rect 92032 2310 92060 2994
rect 92124 2854 92152 36722
rect 96374 36476 96682 36485
rect 96374 36474 96380 36476
rect 96436 36474 96460 36476
rect 96516 36474 96540 36476
rect 96596 36474 96620 36476
rect 96676 36474 96682 36476
rect 96436 36422 96438 36474
rect 96618 36422 96620 36474
rect 96374 36420 96380 36422
rect 96436 36420 96460 36422
rect 96516 36420 96540 36422
rect 96596 36420 96620 36422
rect 96676 36420 96682 36422
rect 96374 36411 96682 36420
rect 96374 35388 96682 35397
rect 96374 35386 96380 35388
rect 96436 35386 96460 35388
rect 96516 35386 96540 35388
rect 96596 35386 96620 35388
rect 96676 35386 96682 35388
rect 96436 35334 96438 35386
rect 96618 35334 96620 35386
rect 96374 35332 96380 35334
rect 96436 35332 96460 35334
rect 96516 35332 96540 35334
rect 96596 35332 96620 35334
rect 96676 35332 96682 35334
rect 96374 35323 96682 35332
rect 96374 34300 96682 34309
rect 96374 34298 96380 34300
rect 96436 34298 96460 34300
rect 96516 34298 96540 34300
rect 96596 34298 96620 34300
rect 96676 34298 96682 34300
rect 96436 34246 96438 34298
rect 96618 34246 96620 34298
rect 96374 34244 96380 34246
rect 96436 34244 96460 34246
rect 96516 34244 96540 34246
rect 96596 34244 96620 34246
rect 96676 34244 96682 34246
rect 96374 34235 96682 34244
rect 92480 33856 92532 33862
rect 92480 33798 92532 33804
rect 92492 3738 92520 33798
rect 96374 33212 96682 33221
rect 96374 33210 96380 33212
rect 96436 33210 96460 33212
rect 96516 33210 96540 33212
rect 96596 33210 96620 33212
rect 96676 33210 96682 33212
rect 96436 33158 96438 33210
rect 96618 33158 96620 33210
rect 96374 33156 96380 33158
rect 96436 33156 96460 33158
rect 96516 33156 96540 33158
rect 96596 33156 96620 33158
rect 96676 33156 96682 33158
rect 96374 33147 96682 33156
rect 96374 32124 96682 32133
rect 96374 32122 96380 32124
rect 96436 32122 96460 32124
rect 96516 32122 96540 32124
rect 96596 32122 96620 32124
rect 96676 32122 96682 32124
rect 96436 32070 96438 32122
rect 96618 32070 96620 32122
rect 96374 32068 96380 32070
rect 96436 32068 96460 32070
rect 96516 32068 96540 32070
rect 96596 32068 96620 32070
rect 96676 32068 96682 32070
rect 96374 32059 96682 32068
rect 96374 31036 96682 31045
rect 96374 31034 96380 31036
rect 96436 31034 96460 31036
rect 96516 31034 96540 31036
rect 96596 31034 96620 31036
rect 96676 31034 96682 31036
rect 96436 30982 96438 31034
rect 96618 30982 96620 31034
rect 96374 30980 96380 30982
rect 96436 30980 96460 30982
rect 96516 30980 96540 30982
rect 96596 30980 96620 30982
rect 96676 30980 96682 30982
rect 96374 30971 96682 30980
rect 96374 29948 96682 29957
rect 96374 29946 96380 29948
rect 96436 29946 96460 29948
rect 96516 29946 96540 29948
rect 96596 29946 96620 29948
rect 96676 29946 96682 29948
rect 96436 29894 96438 29946
rect 96618 29894 96620 29946
rect 96374 29892 96380 29894
rect 96436 29892 96460 29894
rect 96516 29892 96540 29894
rect 96596 29892 96620 29894
rect 96676 29892 96682 29894
rect 96374 29883 96682 29892
rect 96374 28860 96682 28869
rect 96374 28858 96380 28860
rect 96436 28858 96460 28860
rect 96516 28858 96540 28860
rect 96596 28858 96620 28860
rect 96676 28858 96682 28860
rect 96436 28806 96438 28858
rect 96618 28806 96620 28858
rect 96374 28804 96380 28806
rect 96436 28804 96460 28806
rect 96516 28804 96540 28806
rect 96596 28804 96620 28806
rect 96676 28804 96682 28806
rect 96374 28795 96682 28804
rect 96374 27772 96682 27781
rect 96374 27770 96380 27772
rect 96436 27770 96460 27772
rect 96516 27770 96540 27772
rect 96596 27770 96620 27772
rect 96676 27770 96682 27772
rect 96436 27718 96438 27770
rect 96618 27718 96620 27770
rect 96374 27716 96380 27718
rect 96436 27716 96460 27718
rect 96516 27716 96540 27718
rect 96596 27716 96620 27718
rect 96676 27716 96682 27718
rect 96374 27707 96682 27716
rect 96374 26684 96682 26693
rect 96374 26682 96380 26684
rect 96436 26682 96460 26684
rect 96516 26682 96540 26684
rect 96596 26682 96620 26684
rect 96676 26682 96682 26684
rect 96436 26630 96438 26682
rect 96618 26630 96620 26682
rect 96374 26628 96380 26630
rect 96436 26628 96460 26630
rect 96516 26628 96540 26630
rect 96596 26628 96620 26630
rect 96676 26628 96682 26630
rect 96374 26619 96682 26628
rect 96374 25596 96682 25605
rect 96374 25594 96380 25596
rect 96436 25594 96460 25596
rect 96516 25594 96540 25596
rect 96596 25594 96620 25596
rect 96676 25594 96682 25596
rect 96436 25542 96438 25594
rect 96618 25542 96620 25594
rect 96374 25540 96380 25542
rect 96436 25540 96460 25542
rect 96516 25540 96540 25542
rect 96596 25540 96620 25542
rect 96676 25540 96682 25542
rect 96374 25531 96682 25540
rect 96374 24508 96682 24517
rect 96374 24506 96380 24508
rect 96436 24506 96460 24508
rect 96516 24506 96540 24508
rect 96596 24506 96620 24508
rect 96676 24506 96682 24508
rect 96436 24454 96438 24506
rect 96618 24454 96620 24506
rect 96374 24452 96380 24454
rect 96436 24452 96460 24454
rect 96516 24452 96540 24454
rect 96596 24452 96620 24454
rect 96676 24452 96682 24454
rect 96374 24443 96682 24452
rect 96374 23420 96682 23429
rect 96374 23418 96380 23420
rect 96436 23418 96460 23420
rect 96516 23418 96540 23420
rect 96596 23418 96620 23420
rect 96676 23418 96682 23420
rect 96436 23366 96438 23418
rect 96618 23366 96620 23418
rect 96374 23364 96380 23366
rect 96436 23364 96460 23366
rect 96516 23364 96540 23366
rect 96596 23364 96620 23366
rect 96676 23364 96682 23366
rect 96374 23355 96682 23364
rect 96374 22332 96682 22341
rect 96374 22330 96380 22332
rect 96436 22330 96460 22332
rect 96516 22330 96540 22332
rect 96596 22330 96620 22332
rect 96676 22330 96682 22332
rect 96436 22278 96438 22330
rect 96618 22278 96620 22330
rect 96374 22276 96380 22278
rect 96436 22276 96460 22278
rect 96516 22276 96540 22278
rect 96596 22276 96620 22278
rect 96676 22276 96682 22278
rect 96374 22267 96682 22276
rect 96374 21244 96682 21253
rect 96374 21242 96380 21244
rect 96436 21242 96460 21244
rect 96516 21242 96540 21244
rect 96596 21242 96620 21244
rect 96676 21242 96682 21244
rect 96436 21190 96438 21242
rect 96618 21190 96620 21242
rect 96374 21188 96380 21190
rect 96436 21188 96460 21190
rect 96516 21188 96540 21190
rect 96596 21188 96620 21190
rect 96676 21188 96682 21190
rect 96374 21179 96682 21188
rect 96374 20156 96682 20165
rect 96374 20154 96380 20156
rect 96436 20154 96460 20156
rect 96516 20154 96540 20156
rect 96596 20154 96620 20156
rect 96676 20154 96682 20156
rect 96436 20102 96438 20154
rect 96618 20102 96620 20154
rect 96374 20100 96380 20102
rect 96436 20100 96460 20102
rect 96516 20100 96540 20102
rect 96596 20100 96620 20102
rect 96676 20100 96682 20102
rect 96374 20091 96682 20100
rect 96374 19068 96682 19077
rect 96374 19066 96380 19068
rect 96436 19066 96460 19068
rect 96516 19066 96540 19068
rect 96596 19066 96620 19068
rect 96676 19066 96682 19068
rect 96436 19014 96438 19066
rect 96618 19014 96620 19066
rect 96374 19012 96380 19014
rect 96436 19012 96460 19014
rect 96516 19012 96540 19014
rect 96596 19012 96620 19014
rect 96676 19012 96682 19014
rect 96374 19003 96682 19012
rect 96374 17980 96682 17989
rect 96374 17978 96380 17980
rect 96436 17978 96460 17980
rect 96516 17978 96540 17980
rect 96596 17978 96620 17980
rect 96676 17978 96682 17980
rect 96436 17926 96438 17978
rect 96618 17926 96620 17978
rect 96374 17924 96380 17926
rect 96436 17924 96460 17926
rect 96516 17924 96540 17926
rect 96596 17924 96620 17926
rect 96676 17924 96682 17926
rect 96374 17915 96682 17924
rect 96374 16892 96682 16901
rect 96374 16890 96380 16892
rect 96436 16890 96460 16892
rect 96516 16890 96540 16892
rect 96596 16890 96620 16892
rect 96676 16890 96682 16892
rect 96436 16838 96438 16890
rect 96618 16838 96620 16890
rect 96374 16836 96380 16838
rect 96436 16836 96460 16838
rect 96516 16836 96540 16838
rect 96596 16836 96620 16838
rect 96676 16836 96682 16838
rect 96374 16827 96682 16836
rect 96374 15804 96682 15813
rect 96374 15802 96380 15804
rect 96436 15802 96460 15804
rect 96516 15802 96540 15804
rect 96596 15802 96620 15804
rect 96676 15802 96682 15804
rect 96436 15750 96438 15802
rect 96618 15750 96620 15802
rect 96374 15748 96380 15750
rect 96436 15748 96460 15750
rect 96516 15748 96540 15750
rect 96596 15748 96620 15750
rect 96676 15748 96682 15750
rect 96374 15739 96682 15748
rect 96374 14716 96682 14725
rect 96374 14714 96380 14716
rect 96436 14714 96460 14716
rect 96516 14714 96540 14716
rect 96596 14714 96620 14716
rect 96676 14714 96682 14716
rect 96436 14662 96438 14714
rect 96618 14662 96620 14714
rect 96374 14660 96380 14662
rect 96436 14660 96460 14662
rect 96516 14660 96540 14662
rect 96596 14660 96620 14662
rect 96676 14660 96682 14662
rect 96374 14651 96682 14660
rect 96374 13628 96682 13637
rect 96374 13626 96380 13628
rect 96436 13626 96460 13628
rect 96516 13626 96540 13628
rect 96596 13626 96620 13628
rect 96676 13626 96682 13628
rect 96436 13574 96438 13626
rect 96618 13574 96620 13626
rect 96374 13572 96380 13574
rect 96436 13572 96460 13574
rect 96516 13572 96540 13574
rect 96596 13572 96620 13574
rect 96676 13572 96682 13574
rect 96374 13563 96682 13572
rect 96374 12540 96682 12549
rect 96374 12538 96380 12540
rect 96436 12538 96460 12540
rect 96516 12538 96540 12540
rect 96596 12538 96620 12540
rect 96676 12538 96682 12540
rect 96436 12486 96438 12538
rect 96618 12486 96620 12538
rect 96374 12484 96380 12486
rect 96436 12484 96460 12486
rect 96516 12484 96540 12486
rect 96596 12484 96620 12486
rect 96676 12484 96682 12486
rect 96374 12475 96682 12484
rect 96374 11452 96682 11461
rect 96374 11450 96380 11452
rect 96436 11450 96460 11452
rect 96516 11450 96540 11452
rect 96596 11450 96620 11452
rect 96676 11450 96682 11452
rect 96436 11398 96438 11450
rect 96618 11398 96620 11450
rect 96374 11396 96380 11398
rect 96436 11396 96460 11398
rect 96516 11396 96540 11398
rect 96596 11396 96620 11398
rect 96676 11396 96682 11398
rect 96374 11387 96682 11396
rect 96374 10364 96682 10373
rect 96374 10362 96380 10364
rect 96436 10362 96460 10364
rect 96516 10362 96540 10364
rect 96596 10362 96620 10364
rect 96676 10362 96682 10364
rect 96436 10310 96438 10362
rect 96618 10310 96620 10362
rect 96374 10308 96380 10310
rect 96436 10308 96460 10310
rect 96516 10308 96540 10310
rect 96596 10308 96620 10310
rect 96676 10308 96682 10310
rect 96374 10299 96682 10308
rect 96374 9276 96682 9285
rect 96374 9274 96380 9276
rect 96436 9274 96460 9276
rect 96516 9274 96540 9276
rect 96596 9274 96620 9276
rect 96676 9274 96682 9276
rect 96436 9222 96438 9274
rect 96618 9222 96620 9274
rect 96374 9220 96380 9222
rect 96436 9220 96460 9222
rect 96516 9220 96540 9222
rect 96596 9220 96620 9222
rect 96676 9220 96682 9222
rect 96374 9211 96682 9220
rect 96374 8188 96682 8197
rect 96374 8186 96380 8188
rect 96436 8186 96460 8188
rect 96516 8186 96540 8188
rect 96596 8186 96620 8188
rect 96676 8186 96682 8188
rect 96436 8134 96438 8186
rect 96618 8134 96620 8186
rect 96374 8132 96380 8134
rect 96436 8132 96460 8134
rect 96516 8132 96540 8134
rect 96596 8132 96620 8134
rect 96676 8132 96682 8134
rect 96374 8123 96682 8132
rect 96374 7100 96682 7109
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7035 96682 7044
rect 96374 6012 96682 6021
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5947 96682 5956
rect 97632 5364 97684 5370
rect 97632 5306 97684 5312
rect 96804 5228 96856 5234
rect 96804 5170 96856 5176
rect 96988 5228 97040 5234
rect 96988 5170 97040 5176
rect 94044 5160 94096 5166
rect 94044 5102 94096 5108
rect 93952 5024 94004 5030
rect 93952 4966 94004 4972
rect 93964 4622 93992 4966
rect 93952 4616 94004 4622
rect 93952 4558 94004 4564
rect 93860 4072 93912 4078
rect 93860 4014 93912 4020
rect 92480 3732 92532 3738
rect 92480 3674 92532 3680
rect 93872 3126 93900 4014
rect 93964 3602 93992 4558
rect 94056 4554 94084 5102
rect 96632 5098 96752 5114
rect 96620 5092 96752 5098
rect 96672 5086 96752 5092
rect 96620 5034 96672 5040
rect 96374 4924 96682 4933
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4859 96682 4868
rect 94688 4616 94740 4622
rect 94688 4558 94740 4564
rect 94044 4548 94096 4554
rect 94044 4490 94096 4496
rect 94320 4548 94372 4554
rect 94320 4490 94372 4496
rect 94596 4548 94648 4554
rect 94596 4490 94648 4496
rect 93952 3596 94004 3602
rect 93952 3538 94004 3544
rect 93860 3120 93912 3126
rect 93860 3062 93912 3068
rect 94056 3058 94084 4490
rect 94332 4214 94360 4490
rect 94320 4208 94372 4214
rect 94320 4150 94372 4156
rect 94608 4078 94636 4490
rect 94700 4078 94728 4558
rect 96724 4214 96752 5086
rect 96816 4486 96844 5170
rect 97000 4826 97028 5170
rect 96988 4820 97040 4826
rect 96988 4762 97040 4768
rect 97644 4690 97672 5306
rect 100760 5228 100812 5234
rect 100760 5170 100812 5176
rect 100300 5160 100352 5166
rect 100300 5102 100352 5108
rect 100208 5024 100260 5030
rect 100208 4966 100260 4972
rect 97632 4684 97684 4690
rect 97632 4626 97684 4632
rect 100220 4622 100248 4966
rect 100312 4758 100340 5102
rect 100772 4826 100800 5170
rect 100944 5024 100996 5030
rect 100944 4966 100996 4972
rect 100760 4820 100812 4826
rect 100760 4762 100812 4768
rect 100300 4752 100352 4758
rect 100300 4694 100352 4700
rect 100208 4616 100260 4622
rect 100208 4558 100260 4564
rect 96804 4480 96856 4486
rect 96804 4422 96856 4428
rect 99012 4480 99064 4486
rect 99012 4422 99064 4428
rect 96712 4208 96764 4214
rect 96712 4150 96764 4156
rect 97172 4208 97224 4214
rect 97172 4150 97224 4156
rect 94596 4072 94648 4078
rect 94596 4014 94648 4020
rect 94688 4072 94740 4078
rect 94688 4014 94740 4020
rect 94700 3670 94728 4014
rect 96374 3836 96682 3845
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3771 96682 3780
rect 94688 3664 94740 3670
rect 94688 3606 94740 3612
rect 97184 3602 97212 4150
rect 97264 4140 97316 4146
rect 97264 4082 97316 4088
rect 97172 3596 97224 3602
rect 97172 3538 97224 3544
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 94964 3392 95016 3398
rect 94964 3334 95016 3340
rect 94976 3126 95004 3334
rect 95068 3126 95096 3470
rect 97276 3466 97304 4082
rect 98000 3936 98052 3942
rect 98000 3878 98052 3884
rect 98012 3738 98040 3878
rect 98000 3732 98052 3738
rect 98000 3674 98052 3680
rect 97264 3460 97316 3466
rect 97264 3402 97316 3408
rect 96988 3392 97040 3398
rect 96988 3334 97040 3340
rect 94964 3120 95016 3126
rect 94964 3062 95016 3068
rect 95056 3120 95108 3126
rect 95056 3062 95108 3068
rect 94044 3052 94096 3058
rect 94044 2994 94096 3000
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 92112 2848 92164 2854
rect 92112 2790 92164 2796
rect 96252 2848 96304 2854
rect 96252 2790 96304 2796
rect 93952 2508 94004 2514
rect 93952 2450 94004 2456
rect 92388 2440 92440 2446
rect 92388 2382 92440 2388
rect 93400 2440 93452 2446
rect 93400 2382 93452 2388
rect 92400 2310 92428 2382
rect 92020 2304 92072 2310
rect 92020 2246 92072 2252
rect 92388 2304 92440 2310
rect 92388 2246 92440 2252
rect 93136 870 93256 898
rect 93136 800 93164 870
rect 91664 734 91968 762
rect 92294 0 92350 800
rect 93122 0 93178 800
rect 93228 762 93256 870
rect 93412 762 93440 2382
rect 93964 800 93992 2450
rect 95516 2440 95568 2446
rect 95516 2382 95568 2388
rect 95528 800 95556 2382
rect 96264 1306 96292 2790
rect 96374 2748 96682 2757
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2683 96682 2692
rect 96908 2650 96936 2994
rect 97000 2922 97028 3334
rect 98012 2990 98040 3674
rect 98184 3460 98236 3466
rect 98184 3402 98236 3408
rect 98000 2984 98052 2990
rect 98000 2926 98052 2932
rect 96988 2916 97040 2922
rect 96988 2858 97040 2864
rect 98196 2774 98224 3402
rect 98104 2746 98224 2774
rect 96896 2644 96948 2650
rect 96896 2586 96948 2592
rect 98104 2582 98132 2746
rect 98092 2576 98144 2582
rect 98092 2518 98144 2524
rect 99024 2514 99052 4422
rect 100312 3738 100340 4694
rect 100484 4548 100536 4554
rect 100484 4490 100536 4496
rect 100496 4146 100524 4490
rect 100484 4140 100536 4146
rect 100484 4082 100536 4088
rect 100392 4072 100444 4078
rect 100392 4014 100444 4020
rect 100300 3732 100352 3738
rect 100300 3674 100352 3680
rect 100404 3534 100432 4014
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 100392 3528 100444 3534
rect 100392 3470 100444 3476
rect 99300 3346 99328 3470
rect 100772 3398 100800 4762
rect 100956 4622 100984 4966
rect 100944 4616 100996 4622
rect 100944 4558 100996 4564
rect 100956 4282 100984 4558
rect 100944 4276 100996 4282
rect 100944 4218 100996 4224
rect 101128 4276 101180 4282
rect 101128 4218 101180 4224
rect 101140 4146 101168 4218
rect 101312 4208 101364 4214
rect 101312 4150 101364 4156
rect 101128 4140 101180 4146
rect 101128 4082 101180 4088
rect 101324 3602 101352 4150
rect 101784 4146 101812 36790
rect 103796 5364 103848 5370
rect 103796 5306 103848 5312
rect 102324 5160 102376 5166
rect 102324 5102 102376 5108
rect 102336 4486 102364 5102
rect 103808 5030 103836 5306
rect 104532 5228 104584 5234
rect 104532 5170 104584 5176
rect 103796 5024 103848 5030
rect 103796 4966 103848 4972
rect 104544 4826 104572 5170
rect 106464 5160 106516 5166
rect 106464 5102 106516 5108
rect 104532 4820 104584 4826
rect 104532 4762 104584 4768
rect 105084 4752 105136 4758
rect 105084 4694 105136 4700
rect 104716 4616 104768 4622
rect 104716 4558 104768 4564
rect 102324 4480 102376 4486
rect 102324 4422 102376 4428
rect 101496 4140 101548 4146
rect 101496 4082 101548 4088
rect 101772 4140 101824 4146
rect 101772 4082 101824 4088
rect 101312 3596 101364 3602
rect 101312 3538 101364 3544
rect 101508 3534 101536 4082
rect 101680 4072 101732 4078
rect 101680 4014 101732 4020
rect 101692 3602 101720 4014
rect 101784 3602 101812 4082
rect 101680 3596 101732 3602
rect 101680 3538 101732 3544
rect 101772 3596 101824 3602
rect 101772 3538 101824 3544
rect 101496 3528 101548 3534
rect 101496 3470 101548 3476
rect 100760 3392 100812 3398
rect 99300 3318 99420 3346
rect 100760 3334 100812 3340
rect 99012 2508 99064 2514
rect 99012 2450 99064 2456
rect 96712 2440 96764 2446
rect 96712 2382 96764 2388
rect 97908 2440 97960 2446
rect 97908 2382 97960 2388
rect 96724 1834 96752 2382
rect 96712 1828 96764 1834
rect 96712 1770 96764 1776
rect 96264 1278 96384 1306
rect 96356 800 96384 1278
rect 97920 800 97948 2382
rect 99392 1834 99420 3318
rect 99564 3052 99616 3058
rect 99564 2994 99616 3000
rect 100392 3052 100444 3058
rect 100392 2994 100444 3000
rect 99472 2848 99524 2854
rect 99472 2790 99524 2796
rect 99380 1828 99432 1834
rect 99380 1770 99432 1776
rect 99484 800 99512 2790
rect 99576 1698 99604 2994
rect 100300 2576 100352 2582
rect 100300 2518 100352 2524
rect 99564 1692 99616 1698
rect 99564 1634 99616 1640
rect 100312 800 100340 2518
rect 100404 2310 100432 2994
rect 100944 2848 100996 2854
rect 100944 2790 100996 2796
rect 100956 2446 100984 2790
rect 102336 2514 102364 4422
rect 104728 4282 104756 4558
rect 104716 4276 104768 4282
rect 104716 4218 104768 4224
rect 105096 4146 105124 4694
rect 106476 4486 106504 5102
rect 107844 5024 107896 5030
rect 107844 4966 107896 4972
rect 107856 4690 107884 4966
rect 107844 4684 107896 4690
rect 107844 4626 107896 4632
rect 107384 4616 107436 4622
rect 107384 4558 107436 4564
rect 106464 4480 106516 4486
rect 106464 4422 106516 4428
rect 107016 4480 107068 4486
rect 107200 4480 107252 4486
rect 107068 4440 107148 4468
rect 107016 4422 107068 4428
rect 105084 4140 105136 4146
rect 105084 4082 105136 4088
rect 107120 4078 107148 4440
rect 107200 4422 107252 4428
rect 107212 4214 107240 4422
rect 107200 4208 107252 4214
rect 107200 4150 107252 4156
rect 107108 4072 107160 4078
rect 107160 4032 107332 4060
rect 107108 4014 107160 4020
rect 103612 3936 103664 3942
rect 103612 3878 103664 3884
rect 104900 3936 104952 3942
rect 104900 3878 104952 3884
rect 105176 3936 105228 3942
rect 105176 3878 105228 3884
rect 103624 3602 103652 3878
rect 103612 3596 103664 3602
rect 103612 3538 103664 3544
rect 104256 3052 104308 3058
rect 104256 2994 104308 3000
rect 104268 2961 104296 2994
rect 104254 2952 104310 2961
rect 104254 2887 104310 2896
rect 103520 2848 103572 2854
rect 103520 2790 103572 2796
rect 102324 2508 102376 2514
rect 102324 2450 102376 2456
rect 100944 2440 100996 2446
rect 100944 2382 100996 2388
rect 102784 2440 102836 2446
rect 102784 2382 102836 2388
rect 100392 2304 100444 2310
rect 100392 2246 100444 2252
rect 101220 2304 101272 2310
rect 101220 2246 101272 2252
rect 102692 2304 102744 2310
rect 102692 2246 102744 2252
rect 101232 1562 101260 2246
rect 101220 1556 101272 1562
rect 101220 1498 101272 1504
rect 102704 800 102732 2246
rect 102796 1766 102824 2382
rect 102784 1760 102836 1766
rect 102784 1702 102836 1708
rect 103532 800 103560 2790
rect 104912 2446 104940 3878
rect 104992 3052 105044 3058
rect 104992 2994 105044 3000
rect 105004 2650 105032 2994
rect 105188 2922 105216 3878
rect 107304 3097 107332 4032
rect 107396 3738 107424 4558
rect 109696 4010 109724 37198
rect 111734 37020 112042 37029
rect 111734 37018 111740 37020
rect 111796 37018 111820 37020
rect 111876 37018 111900 37020
rect 111956 37018 111980 37020
rect 112036 37018 112042 37020
rect 111796 36966 111798 37018
rect 111978 36966 111980 37018
rect 111734 36964 111740 36966
rect 111796 36964 111820 36966
rect 111876 36964 111900 36966
rect 111956 36964 111980 36966
rect 112036 36964 112042 36966
rect 111734 36955 112042 36964
rect 117240 36922 117268 39199
rect 117884 37126 117912 39200
rect 117504 37120 117556 37126
rect 117504 37062 117556 37068
rect 117872 37120 117924 37126
rect 117872 37062 117924 37068
rect 117228 36916 117280 36922
rect 117228 36858 117280 36864
rect 111734 35932 112042 35941
rect 111734 35930 111740 35932
rect 111796 35930 111820 35932
rect 111876 35930 111900 35932
rect 111956 35930 111980 35932
rect 112036 35930 112042 35932
rect 111796 35878 111798 35930
rect 111978 35878 111980 35930
rect 111734 35876 111740 35878
rect 111796 35876 111820 35878
rect 111876 35876 111900 35878
rect 111956 35876 111980 35878
rect 112036 35876 112042 35878
rect 111734 35867 112042 35876
rect 111734 34844 112042 34853
rect 111734 34842 111740 34844
rect 111796 34842 111820 34844
rect 111876 34842 111900 34844
rect 111956 34842 111980 34844
rect 112036 34842 112042 34844
rect 111796 34790 111798 34842
rect 111978 34790 111980 34842
rect 111734 34788 111740 34790
rect 111796 34788 111820 34790
rect 111876 34788 111900 34790
rect 111956 34788 111980 34790
rect 112036 34788 112042 34790
rect 111734 34779 112042 34788
rect 111734 33756 112042 33765
rect 111734 33754 111740 33756
rect 111796 33754 111820 33756
rect 111876 33754 111900 33756
rect 111956 33754 111980 33756
rect 112036 33754 112042 33756
rect 111796 33702 111798 33754
rect 111978 33702 111980 33754
rect 111734 33700 111740 33702
rect 111796 33700 111820 33702
rect 111876 33700 111900 33702
rect 111956 33700 111980 33702
rect 112036 33700 112042 33702
rect 111734 33691 112042 33700
rect 111734 32668 112042 32677
rect 111734 32666 111740 32668
rect 111796 32666 111820 32668
rect 111876 32666 111900 32668
rect 111956 32666 111980 32668
rect 112036 32666 112042 32668
rect 111796 32614 111798 32666
rect 111978 32614 111980 32666
rect 111734 32612 111740 32614
rect 111796 32612 111820 32614
rect 111876 32612 111900 32614
rect 111956 32612 111980 32614
rect 112036 32612 112042 32614
rect 111734 32603 112042 32612
rect 111734 31580 112042 31589
rect 111734 31578 111740 31580
rect 111796 31578 111820 31580
rect 111876 31578 111900 31580
rect 111956 31578 111980 31580
rect 112036 31578 112042 31580
rect 111796 31526 111798 31578
rect 111978 31526 111980 31578
rect 111734 31524 111740 31526
rect 111796 31524 111820 31526
rect 111876 31524 111900 31526
rect 111956 31524 111980 31526
rect 112036 31524 112042 31526
rect 111734 31515 112042 31524
rect 111734 30492 112042 30501
rect 111734 30490 111740 30492
rect 111796 30490 111820 30492
rect 111876 30490 111900 30492
rect 111956 30490 111980 30492
rect 112036 30490 112042 30492
rect 111796 30438 111798 30490
rect 111978 30438 111980 30490
rect 111734 30436 111740 30438
rect 111796 30436 111820 30438
rect 111876 30436 111900 30438
rect 111956 30436 111980 30438
rect 112036 30436 112042 30438
rect 111734 30427 112042 30436
rect 112444 29504 112496 29510
rect 112444 29446 112496 29452
rect 111734 29404 112042 29413
rect 111734 29402 111740 29404
rect 111796 29402 111820 29404
rect 111876 29402 111900 29404
rect 111956 29402 111980 29404
rect 112036 29402 112042 29404
rect 111796 29350 111798 29402
rect 111978 29350 111980 29402
rect 111734 29348 111740 29350
rect 111796 29348 111820 29350
rect 111876 29348 111900 29350
rect 111956 29348 111980 29350
rect 112036 29348 112042 29350
rect 111734 29339 112042 29348
rect 111734 28316 112042 28325
rect 111734 28314 111740 28316
rect 111796 28314 111820 28316
rect 111876 28314 111900 28316
rect 111956 28314 111980 28316
rect 112036 28314 112042 28316
rect 111796 28262 111798 28314
rect 111978 28262 111980 28314
rect 111734 28260 111740 28262
rect 111796 28260 111820 28262
rect 111876 28260 111900 28262
rect 111956 28260 111980 28262
rect 112036 28260 112042 28262
rect 111734 28251 112042 28260
rect 111734 27228 112042 27237
rect 111734 27226 111740 27228
rect 111796 27226 111820 27228
rect 111876 27226 111900 27228
rect 111956 27226 111980 27228
rect 112036 27226 112042 27228
rect 111796 27174 111798 27226
rect 111978 27174 111980 27226
rect 111734 27172 111740 27174
rect 111796 27172 111820 27174
rect 111876 27172 111900 27174
rect 111956 27172 111980 27174
rect 112036 27172 112042 27174
rect 111734 27163 112042 27172
rect 111734 26140 112042 26149
rect 111734 26138 111740 26140
rect 111796 26138 111820 26140
rect 111876 26138 111900 26140
rect 111956 26138 111980 26140
rect 112036 26138 112042 26140
rect 111796 26086 111798 26138
rect 111978 26086 111980 26138
rect 111734 26084 111740 26086
rect 111796 26084 111820 26086
rect 111876 26084 111900 26086
rect 111956 26084 111980 26086
rect 112036 26084 112042 26086
rect 111734 26075 112042 26084
rect 111734 25052 112042 25061
rect 111734 25050 111740 25052
rect 111796 25050 111820 25052
rect 111876 25050 111900 25052
rect 111956 25050 111980 25052
rect 112036 25050 112042 25052
rect 111796 24998 111798 25050
rect 111978 24998 111980 25050
rect 111734 24996 111740 24998
rect 111796 24996 111820 24998
rect 111876 24996 111900 24998
rect 111956 24996 111980 24998
rect 112036 24996 112042 24998
rect 111734 24987 112042 24996
rect 111734 23964 112042 23973
rect 111734 23962 111740 23964
rect 111796 23962 111820 23964
rect 111876 23962 111900 23964
rect 111956 23962 111980 23964
rect 112036 23962 112042 23964
rect 111796 23910 111798 23962
rect 111978 23910 111980 23962
rect 111734 23908 111740 23910
rect 111796 23908 111820 23910
rect 111876 23908 111900 23910
rect 111956 23908 111980 23910
rect 112036 23908 112042 23910
rect 111734 23899 112042 23908
rect 111734 22876 112042 22885
rect 111734 22874 111740 22876
rect 111796 22874 111820 22876
rect 111876 22874 111900 22876
rect 111956 22874 111980 22876
rect 112036 22874 112042 22876
rect 111796 22822 111798 22874
rect 111978 22822 111980 22874
rect 111734 22820 111740 22822
rect 111796 22820 111820 22822
rect 111876 22820 111900 22822
rect 111956 22820 111980 22822
rect 112036 22820 112042 22822
rect 111734 22811 112042 22820
rect 111734 21788 112042 21797
rect 111734 21786 111740 21788
rect 111796 21786 111820 21788
rect 111876 21786 111900 21788
rect 111956 21786 111980 21788
rect 112036 21786 112042 21788
rect 111796 21734 111798 21786
rect 111978 21734 111980 21786
rect 111734 21732 111740 21734
rect 111796 21732 111820 21734
rect 111876 21732 111900 21734
rect 111956 21732 111980 21734
rect 112036 21732 112042 21734
rect 111734 21723 112042 21732
rect 111734 20700 112042 20709
rect 111734 20698 111740 20700
rect 111796 20698 111820 20700
rect 111876 20698 111900 20700
rect 111956 20698 111980 20700
rect 112036 20698 112042 20700
rect 111796 20646 111798 20698
rect 111978 20646 111980 20698
rect 111734 20644 111740 20646
rect 111796 20644 111820 20646
rect 111876 20644 111900 20646
rect 111956 20644 111980 20646
rect 112036 20644 112042 20646
rect 111734 20635 112042 20644
rect 111734 19612 112042 19621
rect 111734 19610 111740 19612
rect 111796 19610 111820 19612
rect 111876 19610 111900 19612
rect 111956 19610 111980 19612
rect 112036 19610 112042 19612
rect 111796 19558 111798 19610
rect 111978 19558 111980 19610
rect 111734 19556 111740 19558
rect 111796 19556 111820 19558
rect 111876 19556 111900 19558
rect 111956 19556 111980 19558
rect 112036 19556 112042 19558
rect 111734 19547 112042 19556
rect 111734 18524 112042 18533
rect 111734 18522 111740 18524
rect 111796 18522 111820 18524
rect 111876 18522 111900 18524
rect 111956 18522 111980 18524
rect 112036 18522 112042 18524
rect 111796 18470 111798 18522
rect 111978 18470 111980 18522
rect 111734 18468 111740 18470
rect 111796 18468 111820 18470
rect 111876 18468 111900 18470
rect 111956 18468 111980 18470
rect 112036 18468 112042 18470
rect 111734 18459 112042 18468
rect 111734 17436 112042 17445
rect 111734 17434 111740 17436
rect 111796 17434 111820 17436
rect 111876 17434 111900 17436
rect 111956 17434 111980 17436
rect 112036 17434 112042 17436
rect 111796 17382 111798 17434
rect 111978 17382 111980 17434
rect 111734 17380 111740 17382
rect 111796 17380 111820 17382
rect 111876 17380 111900 17382
rect 111956 17380 111980 17382
rect 112036 17380 112042 17382
rect 111734 17371 112042 17380
rect 111734 16348 112042 16357
rect 111734 16346 111740 16348
rect 111796 16346 111820 16348
rect 111876 16346 111900 16348
rect 111956 16346 111980 16348
rect 112036 16346 112042 16348
rect 111796 16294 111798 16346
rect 111978 16294 111980 16346
rect 111734 16292 111740 16294
rect 111796 16292 111820 16294
rect 111876 16292 111900 16294
rect 111956 16292 111980 16294
rect 112036 16292 112042 16294
rect 111734 16283 112042 16292
rect 111734 15260 112042 15269
rect 111734 15258 111740 15260
rect 111796 15258 111820 15260
rect 111876 15258 111900 15260
rect 111956 15258 111980 15260
rect 112036 15258 112042 15260
rect 111796 15206 111798 15258
rect 111978 15206 111980 15258
rect 111734 15204 111740 15206
rect 111796 15204 111820 15206
rect 111876 15204 111900 15206
rect 111956 15204 111980 15206
rect 112036 15204 112042 15206
rect 111734 15195 112042 15204
rect 111734 14172 112042 14181
rect 111734 14170 111740 14172
rect 111796 14170 111820 14172
rect 111876 14170 111900 14172
rect 111956 14170 111980 14172
rect 112036 14170 112042 14172
rect 111796 14118 111798 14170
rect 111978 14118 111980 14170
rect 111734 14116 111740 14118
rect 111796 14116 111820 14118
rect 111876 14116 111900 14118
rect 111956 14116 111980 14118
rect 112036 14116 112042 14118
rect 111734 14107 112042 14116
rect 111734 13084 112042 13093
rect 111734 13082 111740 13084
rect 111796 13082 111820 13084
rect 111876 13082 111900 13084
rect 111956 13082 111980 13084
rect 112036 13082 112042 13084
rect 111796 13030 111798 13082
rect 111978 13030 111980 13082
rect 111734 13028 111740 13030
rect 111796 13028 111820 13030
rect 111876 13028 111900 13030
rect 111956 13028 111980 13030
rect 112036 13028 112042 13030
rect 111734 13019 112042 13028
rect 111734 11996 112042 12005
rect 111734 11994 111740 11996
rect 111796 11994 111820 11996
rect 111876 11994 111900 11996
rect 111956 11994 111980 11996
rect 112036 11994 112042 11996
rect 111796 11942 111798 11994
rect 111978 11942 111980 11994
rect 111734 11940 111740 11942
rect 111796 11940 111820 11942
rect 111876 11940 111900 11942
rect 111956 11940 111980 11942
rect 112036 11940 112042 11942
rect 111734 11931 112042 11940
rect 111734 10908 112042 10917
rect 111734 10906 111740 10908
rect 111796 10906 111820 10908
rect 111876 10906 111900 10908
rect 111956 10906 111980 10908
rect 112036 10906 112042 10908
rect 111796 10854 111798 10906
rect 111978 10854 111980 10906
rect 111734 10852 111740 10854
rect 111796 10852 111820 10854
rect 111876 10852 111900 10854
rect 111956 10852 111980 10854
rect 112036 10852 112042 10854
rect 111734 10843 112042 10852
rect 111734 9820 112042 9829
rect 111734 9818 111740 9820
rect 111796 9818 111820 9820
rect 111876 9818 111900 9820
rect 111956 9818 111980 9820
rect 112036 9818 112042 9820
rect 111796 9766 111798 9818
rect 111978 9766 111980 9818
rect 111734 9764 111740 9766
rect 111796 9764 111820 9766
rect 111876 9764 111900 9766
rect 111956 9764 111980 9766
rect 112036 9764 112042 9766
rect 111734 9755 112042 9764
rect 111734 8732 112042 8741
rect 111734 8730 111740 8732
rect 111796 8730 111820 8732
rect 111876 8730 111900 8732
rect 111956 8730 111980 8732
rect 112036 8730 112042 8732
rect 111796 8678 111798 8730
rect 111978 8678 111980 8730
rect 111734 8676 111740 8678
rect 111796 8676 111820 8678
rect 111876 8676 111900 8678
rect 111956 8676 111980 8678
rect 112036 8676 112042 8678
rect 111734 8667 112042 8676
rect 111734 7644 112042 7653
rect 111734 7642 111740 7644
rect 111796 7642 111820 7644
rect 111876 7642 111900 7644
rect 111956 7642 111980 7644
rect 112036 7642 112042 7644
rect 111796 7590 111798 7642
rect 111978 7590 111980 7642
rect 111734 7588 111740 7590
rect 111796 7588 111820 7590
rect 111876 7588 111900 7590
rect 111956 7588 111980 7590
rect 112036 7588 112042 7590
rect 111734 7579 112042 7588
rect 111734 6556 112042 6565
rect 111734 6554 111740 6556
rect 111796 6554 111820 6556
rect 111876 6554 111900 6556
rect 111956 6554 111980 6556
rect 112036 6554 112042 6556
rect 111796 6502 111798 6554
rect 111978 6502 111980 6554
rect 111734 6500 111740 6502
rect 111796 6500 111820 6502
rect 111876 6500 111900 6502
rect 111956 6500 111980 6502
rect 112036 6500 112042 6502
rect 111734 6491 112042 6500
rect 111734 5468 112042 5477
rect 111734 5466 111740 5468
rect 111796 5466 111820 5468
rect 111876 5466 111900 5468
rect 111956 5466 111980 5468
rect 112036 5466 112042 5468
rect 111796 5414 111798 5466
rect 111978 5414 111980 5466
rect 111734 5412 111740 5414
rect 111796 5412 111820 5414
rect 111876 5412 111900 5414
rect 111956 5412 111980 5414
rect 112036 5412 112042 5414
rect 111734 5403 112042 5412
rect 109960 4752 110012 4758
rect 109960 4694 110012 4700
rect 109684 4004 109736 4010
rect 109684 3946 109736 3952
rect 108488 3936 108540 3942
rect 108488 3878 108540 3884
rect 107384 3732 107436 3738
rect 107384 3674 107436 3680
rect 108500 3602 108528 3878
rect 109776 3732 109828 3738
rect 109776 3674 109828 3680
rect 108488 3596 108540 3602
rect 108488 3538 108540 3544
rect 108396 3528 108448 3534
rect 108396 3470 108448 3476
rect 107290 3088 107346 3097
rect 107290 3023 107292 3032
rect 107344 3023 107346 3032
rect 108304 3052 108356 3058
rect 107292 2994 107344 3000
rect 108304 2994 108356 3000
rect 105176 2916 105228 2922
rect 105176 2858 105228 2864
rect 105084 2848 105136 2854
rect 105084 2790 105136 2796
rect 104992 2644 105044 2650
rect 104992 2586 105044 2592
rect 104900 2440 104952 2446
rect 104900 2382 104952 2388
rect 105096 800 105124 2790
rect 108316 2650 108344 2994
rect 108304 2644 108356 2650
rect 108304 2586 108356 2592
rect 107568 2440 107620 2446
rect 107568 2382 107620 2388
rect 107476 2304 107528 2310
rect 107476 2246 107528 2252
rect 107488 800 107516 2246
rect 107580 2106 107608 2382
rect 107568 2100 107620 2106
rect 107568 2042 107620 2048
rect 108408 1850 108436 3470
rect 109788 2922 109816 3674
rect 109776 2916 109828 2922
rect 109776 2858 109828 2864
rect 109788 2446 109816 2858
rect 109972 2854 110000 4694
rect 112456 4690 112484 29446
rect 117226 12200 117282 12209
rect 117226 12135 117228 12144
rect 117280 12135 117282 12144
rect 117228 12106 117280 12112
rect 114468 6656 114520 6662
rect 114468 6598 114520 6604
rect 114480 5098 114508 6598
rect 114468 5092 114520 5098
rect 114468 5034 114520 5040
rect 112444 4684 112496 4690
rect 112444 4626 112496 4632
rect 111156 4480 111208 4486
rect 111156 4422 111208 4428
rect 112352 4480 112404 4486
rect 112352 4422 112404 4428
rect 111168 4214 111196 4422
rect 111734 4380 112042 4389
rect 111734 4378 111740 4380
rect 111796 4378 111820 4380
rect 111876 4378 111900 4380
rect 111956 4378 111980 4380
rect 112036 4378 112042 4380
rect 111796 4326 111798 4378
rect 111978 4326 111980 4378
rect 111734 4324 111740 4326
rect 111796 4324 111820 4326
rect 111876 4324 111900 4326
rect 111956 4324 111980 4326
rect 112036 4324 112042 4326
rect 111734 4315 112042 4324
rect 112364 4282 112392 4422
rect 112352 4276 112404 4282
rect 112352 4218 112404 4224
rect 111156 4208 111208 4214
rect 111156 4150 111208 4156
rect 110972 3936 111024 3942
rect 110972 3878 111024 3884
rect 110984 3097 111012 3878
rect 111996 3466 112116 3482
rect 112364 3466 112392 4218
rect 117516 3738 117544 37062
rect 118054 35048 118110 35057
rect 118054 34983 118110 34992
rect 118068 34950 118096 34983
rect 118056 34944 118108 34950
rect 118056 34886 118108 34892
rect 118056 33856 118108 33862
rect 118056 33798 118108 33804
rect 118068 33561 118096 33798
rect 118054 33552 118110 33561
rect 118054 33487 118110 33496
rect 117964 29572 118016 29578
rect 117964 29514 118016 29520
rect 117976 29345 118004 29514
rect 117962 29336 118018 29345
rect 117962 29271 118018 29280
rect 118056 26784 118108 26790
rect 118056 26726 118108 26732
rect 118068 26489 118096 26726
rect 118054 26480 118110 26489
rect 118054 26415 118110 26424
rect 118054 23624 118110 23633
rect 118054 23559 118056 23568
rect 118108 23559 118110 23568
rect 118056 23530 118108 23536
rect 118056 22432 118108 22438
rect 118056 22374 118108 22380
rect 118068 22137 118096 22374
rect 118054 22128 118110 22137
rect 118054 22063 118110 22072
rect 117780 20868 117832 20874
rect 117780 20810 117832 20816
rect 117792 20777 117820 20810
rect 117778 20768 117834 20777
rect 117778 20703 117834 20712
rect 118056 19508 118108 19514
rect 118056 19450 118108 19456
rect 117872 19372 117924 19378
rect 117872 19314 117924 19320
rect 117884 18630 117912 19314
rect 118068 19281 118096 19450
rect 118054 19272 118110 19281
rect 118054 19207 118110 19216
rect 117872 18624 117924 18630
rect 117872 18566 117924 18572
rect 117780 18284 117832 18290
rect 117780 18226 117832 18232
rect 117792 17921 117820 18226
rect 117872 18080 117924 18086
rect 117872 18022 117924 18028
rect 117778 17912 117834 17921
rect 117778 17847 117834 17856
rect 117780 15428 117832 15434
rect 117780 15370 117832 15376
rect 117792 15065 117820 15370
rect 117778 15056 117834 15065
rect 117778 14991 117834 15000
rect 117884 6914 117912 18022
rect 117792 6886 117912 6914
rect 117792 5302 117820 6886
rect 117964 6724 118016 6730
rect 117964 6666 118016 6672
rect 117976 6497 118004 6666
rect 117962 6488 118018 6497
rect 117962 6423 118018 6432
rect 117780 5296 117832 5302
rect 117780 5238 117832 5244
rect 118056 5024 118108 5030
rect 118054 4992 118056 5001
rect 118108 4992 118110 5001
rect 118054 4927 118110 4936
rect 117964 4208 118016 4214
rect 117964 4150 118016 4156
rect 117504 3732 117556 3738
rect 117504 3674 117556 3680
rect 117976 3641 118004 4150
rect 117962 3632 118018 3641
rect 117962 3567 118018 3576
rect 115572 3528 115624 3534
rect 115572 3470 115624 3476
rect 117412 3528 117464 3534
rect 117412 3470 117464 3476
rect 111984 3460 112116 3466
rect 112036 3454 112116 3460
rect 111984 3402 112036 3408
rect 111734 3292 112042 3301
rect 111734 3290 111740 3292
rect 111796 3290 111820 3292
rect 111876 3290 111900 3292
rect 111956 3290 111980 3292
rect 112036 3290 112042 3292
rect 111796 3238 111798 3290
rect 111978 3238 111980 3290
rect 111734 3236 111740 3238
rect 111796 3236 111820 3238
rect 111876 3236 111900 3238
rect 111956 3236 111980 3238
rect 112036 3236 112042 3238
rect 111734 3227 112042 3236
rect 110970 3088 111026 3097
rect 110970 3023 111026 3032
rect 111432 3052 111484 3058
rect 110984 2990 111012 3023
rect 111432 2994 111484 3000
rect 110972 2984 111024 2990
rect 110972 2926 111024 2932
rect 109960 2848 110012 2854
rect 109960 2790 110012 2796
rect 109972 2514 110000 2790
rect 109960 2508 110012 2514
rect 109960 2450 110012 2456
rect 109776 2440 109828 2446
rect 109776 2382 109828 2388
rect 109868 2440 109920 2446
rect 109868 2382 109920 2388
rect 108316 1822 108436 1850
rect 108316 800 108344 1822
rect 109880 800 109908 2382
rect 110696 2372 110748 2378
rect 110696 2314 110748 2320
rect 110708 800 110736 2314
rect 111444 1034 111472 2994
rect 112088 2802 112116 3454
rect 112352 3460 112404 3466
rect 112352 3402 112404 3408
rect 112628 3392 112680 3398
rect 112628 3334 112680 3340
rect 112640 3194 112668 3334
rect 115584 3194 115612 3470
rect 112628 3188 112680 3194
rect 112628 3130 112680 3136
rect 115572 3188 115624 3194
rect 115572 3130 115624 3136
rect 112260 3052 112312 3058
rect 112260 2994 112312 3000
rect 114836 3052 114888 3058
rect 114836 2994 114888 3000
rect 112168 2848 112220 2854
rect 112088 2796 112168 2802
rect 112088 2790 112220 2796
rect 112088 2774 112208 2790
rect 112088 2446 112116 2774
rect 112272 2650 112300 2994
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 112260 2644 112312 2650
rect 112260 2586 112312 2592
rect 112352 2576 112404 2582
rect 112352 2518 112404 2524
rect 112076 2440 112128 2446
rect 112076 2382 112128 2388
rect 111734 2204 112042 2213
rect 111734 2202 111740 2204
rect 111796 2202 111820 2204
rect 111876 2202 111900 2204
rect 111956 2202 111980 2204
rect 112036 2202 112042 2204
rect 111796 2150 111798 2202
rect 111978 2150 111980 2202
rect 111734 2148 111740 2150
rect 111796 2148 111820 2150
rect 111876 2148 111900 2150
rect 111956 2148 111980 2150
rect 112036 2148 112042 2150
rect 111734 2139 112042 2148
rect 111444 1006 111564 1034
rect 111536 800 111564 1006
rect 112364 800 112392 2518
rect 112812 2440 112864 2446
rect 112812 2382 112864 2388
rect 114560 2440 114612 2446
rect 114560 2382 114612 2388
rect 112824 2310 112852 2382
rect 112812 2304 112864 2310
rect 112812 2246 112864 2252
rect 113916 2304 113968 2310
rect 113916 2246 113968 2252
rect 112824 1494 112852 2246
rect 112812 1488 112864 1494
rect 112812 1430 112864 1436
rect 113928 800 113956 2246
rect 114572 2038 114600 2382
rect 114560 2032 114612 2038
rect 114560 1974 114612 1980
rect 114756 800 114784 2790
rect 114848 1630 114876 2994
rect 115480 2440 115532 2446
rect 115480 2382 115532 2388
rect 115848 2440 115900 2446
rect 115848 2382 115900 2388
rect 117136 2440 117188 2446
rect 117136 2382 117188 2388
rect 117228 2440 117280 2446
rect 117228 2382 117280 2388
rect 114836 1624 114888 1630
rect 114836 1566 114888 1572
rect 115492 800 115520 2382
rect 115860 1834 115888 2382
rect 116308 2304 116360 2310
rect 116308 2246 116360 2252
rect 115848 1828 115900 1834
rect 115848 1770 115900 1776
rect 116320 800 116348 2246
rect 117148 1902 117176 2382
rect 117240 1970 117268 2382
rect 117424 2378 117452 3470
rect 118148 3392 118200 3398
rect 118148 3334 118200 3340
rect 117964 3052 118016 3058
rect 117964 2994 118016 3000
rect 117412 2372 117464 2378
rect 117412 2314 117464 2320
rect 117872 2304 117924 2310
rect 117872 2246 117924 2252
rect 117228 1964 117280 1970
rect 117228 1906 117280 1912
rect 117136 1896 117188 1902
rect 117136 1838 117188 1844
rect 117884 800 117912 2246
rect 117976 2145 118004 2994
rect 117962 2136 118018 2145
rect 117962 2071 118018 2080
rect 93228 734 93440 762
rect 93950 0 94006 800
rect 94686 0 94742 800
rect 95514 0 95570 800
rect 96342 0 96398 800
rect 97078 0 97134 800
rect 97906 0 97962 800
rect 98734 0 98790 800
rect 99470 0 99526 800
rect 100298 0 100354 800
rect 101126 0 101182 800
rect 101954 0 102010 800
rect 102690 0 102746 800
rect 103518 0 103574 800
rect 104346 0 104402 800
rect 105082 0 105138 800
rect 105910 0 105966 800
rect 106738 0 106794 800
rect 107474 0 107530 800
rect 108302 0 108358 800
rect 109130 0 109186 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115478 0 115534 800
rect 116306 0 116362 800
rect 117134 0 117190 800
rect 117870 0 117926 800
rect 118160 785 118188 3334
rect 118146 776 118202 785
rect 118146 711 118202 720
rect 118698 0 118754 800
rect 119526 0 119582 800
<< via2 >>
rect 1582 37460 1638 37496
rect 2778 39072 2834 39128
rect 1582 37440 1584 37460
rect 1584 37440 1636 37460
rect 1636 37440 1638 37460
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 117226 39208 117282 39264
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 1490 35808 1546 35864
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 1582 34176 1638 34232
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 1398 25744 1454 25800
rect 1398 22480 1454 22536
rect 1398 19080 1454 19136
rect 1398 17448 1454 17504
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 1582 32408 1638 32464
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 1582 29144 1638 29200
rect 1582 24112 1638 24168
rect 1582 9152 1638 9208
rect 1582 7520 1638 7576
rect 1858 14184 1914 14240
rect 1858 10784 1914 10840
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1398 856 1454 912
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 39670 2932 39672 2952
rect 39672 2932 39724 2952
rect 39724 2932 39726 2952
rect 39670 2896 39726 2932
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 47582 2932 47584 2952
rect 47584 2932 47636 2952
rect 47636 2932 47638 2952
rect 47582 2896 47638 2932
rect 50618 2896 50674 2952
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 81020 37018 81076 37020
rect 81100 37018 81156 37020
rect 81180 37018 81236 37020
rect 81260 37018 81316 37020
rect 81020 36966 81066 37018
rect 81066 36966 81076 37018
rect 81100 36966 81130 37018
rect 81130 36966 81142 37018
rect 81142 36966 81156 37018
rect 81180 36966 81194 37018
rect 81194 36966 81206 37018
rect 81206 36966 81236 37018
rect 81260 36966 81270 37018
rect 81270 36966 81316 37018
rect 81020 36964 81076 36966
rect 81100 36964 81156 36966
rect 81180 36964 81236 36966
rect 81260 36964 81316 36966
rect 81020 35930 81076 35932
rect 81100 35930 81156 35932
rect 81180 35930 81236 35932
rect 81260 35930 81316 35932
rect 81020 35878 81066 35930
rect 81066 35878 81076 35930
rect 81100 35878 81130 35930
rect 81130 35878 81142 35930
rect 81142 35878 81156 35930
rect 81180 35878 81194 35930
rect 81194 35878 81206 35930
rect 81206 35878 81236 35930
rect 81260 35878 81270 35930
rect 81270 35878 81316 35930
rect 81020 35876 81076 35878
rect 81100 35876 81156 35878
rect 81180 35876 81236 35878
rect 81260 35876 81316 35878
rect 81020 34842 81076 34844
rect 81100 34842 81156 34844
rect 81180 34842 81236 34844
rect 81260 34842 81316 34844
rect 81020 34790 81066 34842
rect 81066 34790 81076 34842
rect 81100 34790 81130 34842
rect 81130 34790 81142 34842
rect 81142 34790 81156 34842
rect 81180 34790 81194 34842
rect 81194 34790 81206 34842
rect 81206 34790 81236 34842
rect 81260 34790 81270 34842
rect 81270 34790 81316 34842
rect 81020 34788 81076 34790
rect 81100 34788 81156 34790
rect 81180 34788 81236 34790
rect 81260 34788 81316 34790
rect 81020 33754 81076 33756
rect 81100 33754 81156 33756
rect 81180 33754 81236 33756
rect 81260 33754 81316 33756
rect 81020 33702 81066 33754
rect 81066 33702 81076 33754
rect 81100 33702 81130 33754
rect 81130 33702 81142 33754
rect 81142 33702 81156 33754
rect 81180 33702 81194 33754
rect 81194 33702 81206 33754
rect 81206 33702 81236 33754
rect 81260 33702 81270 33754
rect 81270 33702 81316 33754
rect 81020 33700 81076 33702
rect 81100 33700 81156 33702
rect 81180 33700 81236 33702
rect 81260 33700 81316 33702
rect 81020 32666 81076 32668
rect 81100 32666 81156 32668
rect 81180 32666 81236 32668
rect 81260 32666 81316 32668
rect 81020 32614 81066 32666
rect 81066 32614 81076 32666
rect 81100 32614 81130 32666
rect 81130 32614 81142 32666
rect 81142 32614 81156 32666
rect 81180 32614 81194 32666
rect 81194 32614 81206 32666
rect 81206 32614 81236 32666
rect 81260 32614 81270 32666
rect 81270 32614 81316 32666
rect 81020 32612 81076 32614
rect 81100 32612 81156 32614
rect 81180 32612 81236 32614
rect 81260 32612 81316 32614
rect 81020 31578 81076 31580
rect 81100 31578 81156 31580
rect 81180 31578 81236 31580
rect 81260 31578 81316 31580
rect 81020 31526 81066 31578
rect 81066 31526 81076 31578
rect 81100 31526 81130 31578
rect 81130 31526 81142 31578
rect 81142 31526 81156 31578
rect 81180 31526 81194 31578
rect 81194 31526 81206 31578
rect 81206 31526 81236 31578
rect 81260 31526 81270 31578
rect 81270 31526 81316 31578
rect 81020 31524 81076 31526
rect 81100 31524 81156 31526
rect 81180 31524 81236 31526
rect 81260 31524 81316 31526
rect 81020 30490 81076 30492
rect 81100 30490 81156 30492
rect 81180 30490 81236 30492
rect 81260 30490 81316 30492
rect 81020 30438 81066 30490
rect 81066 30438 81076 30490
rect 81100 30438 81130 30490
rect 81130 30438 81142 30490
rect 81142 30438 81156 30490
rect 81180 30438 81194 30490
rect 81194 30438 81206 30490
rect 81206 30438 81236 30490
rect 81260 30438 81270 30490
rect 81270 30438 81316 30490
rect 81020 30436 81076 30438
rect 81100 30436 81156 30438
rect 81180 30436 81236 30438
rect 81260 30436 81316 30438
rect 81020 29402 81076 29404
rect 81100 29402 81156 29404
rect 81180 29402 81236 29404
rect 81260 29402 81316 29404
rect 81020 29350 81066 29402
rect 81066 29350 81076 29402
rect 81100 29350 81130 29402
rect 81130 29350 81142 29402
rect 81142 29350 81156 29402
rect 81180 29350 81194 29402
rect 81194 29350 81206 29402
rect 81206 29350 81236 29402
rect 81260 29350 81270 29402
rect 81270 29350 81316 29402
rect 81020 29348 81076 29350
rect 81100 29348 81156 29350
rect 81180 29348 81236 29350
rect 81260 29348 81316 29350
rect 81020 28314 81076 28316
rect 81100 28314 81156 28316
rect 81180 28314 81236 28316
rect 81260 28314 81316 28316
rect 81020 28262 81066 28314
rect 81066 28262 81076 28314
rect 81100 28262 81130 28314
rect 81130 28262 81142 28314
rect 81142 28262 81156 28314
rect 81180 28262 81194 28314
rect 81194 28262 81206 28314
rect 81206 28262 81236 28314
rect 81260 28262 81270 28314
rect 81270 28262 81316 28314
rect 81020 28260 81076 28262
rect 81100 28260 81156 28262
rect 81180 28260 81236 28262
rect 81260 28260 81316 28262
rect 81020 27226 81076 27228
rect 81100 27226 81156 27228
rect 81180 27226 81236 27228
rect 81260 27226 81316 27228
rect 81020 27174 81066 27226
rect 81066 27174 81076 27226
rect 81100 27174 81130 27226
rect 81130 27174 81142 27226
rect 81142 27174 81156 27226
rect 81180 27174 81194 27226
rect 81194 27174 81206 27226
rect 81206 27174 81236 27226
rect 81260 27174 81270 27226
rect 81270 27174 81316 27226
rect 81020 27172 81076 27174
rect 81100 27172 81156 27174
rect 81180 27172 81236 27174
rect 81260 27172 81316 27174
rect 81020 26138 81076 26140
rect 81100 26138 81156 26140
rect 81180 26138 81236 26140
rect 81260 26138 81316 26140
rect 81020 26086 81066 26138
rect 81066 26086 81076 26138
rect 81100 26086 81130 26138
rect 81130 26086 81142 26138
rect 81142 26086 81156 26138
rect 81180 26086 81194 26138
rect 81194 26086 81206 26138
rect 81206 26086 81236 26138
rect 81260 26086 81270 26138
rect 81270 26086 81316 26138
rect 81020 26084 81076 26086
rect 81100 26084 81156 26086
rect 81180 26084 81236 26086
rect 81260 26084 81316 26086
rect 81020 25050 81076 25052
rect 81100 25050 81156 25052
rect 81180 25050 81236 25052
rect 81260 25050 81316 25052
rect 81020 24998 81066 25050
rect 81066 24998 81076 25050
rect 81100 24998 81130 25050
rect 81130 24998 81142 25050
rect 81142 24998 81156 25050
rect 81180 24998 81194 25050
rect 81194 24998 81206 25050
rect 81206 24998 81236 25050
rect 81260 24998 81270 25050
rect 81270 24998 81316 25050
rect 81020 24996 81076 24998
rect 81100 24996 81156 24998
rect 81180 24996 81236 24998
rect 81260 24996 81316 24998
rect 81020 23962 81076 23964
rect 81100 23962 81156 23964
rect 81180 23962 81236 23964
rect 81260 23962 81316 23964
rect 81020 23910 81066 23962
rect 81066 23910 81076 23962
rect 81100 23910 81130 23962
rect 81130 23910 81142 23962
rect 81142 23910 81156 23962
rect 81180 23910 81194 23962
rect 81194 23910 81206 23962
rect 81206 23910 81236 23962
rect 81260 23910 81270 23962
rect 81270 23910 81316 23962
rect 81020 23908 81076 23910
rect 81100 23908 81156 23910
rect 81180 23908 81236 23910
rect 81260 23908 81316 23910
rect 81020 22874 81076 22876
rect 81100 22874 81156 22876
rect 81180 22874 81236 22876
rect 81260 22874 81316 22876
rect 81020 22822 81066 22874
rect 81066 22822 81076 22874
rect 81100 22822 81130 22874
rect 81130 22822 81142 22874
rect 81142 22822 81156 22874
rect 81180 22822 81194 22874
rect 81194 22822 81206 22874
rect 81206 22822 81236 22874
rect 81260 22822 81270 22874
rect 81270 22822 81316 22874
rect 81020 22820 81076 22822
rect 81100 22820 81156 22822
rect 81180 22820 81236 22822
rect 81260 22820 81316 22822
rect 81020 21786 81076 21788
rect 81100 21786 81156 21788
rect 81180 21786 81236 21788
rect 81260 21786 81316 21788
rect 81020 21734 81066 21786
rect 81066 21734 81076 21786
rect 81100 21734 81130 21786
rect 81130 21734 81142 21786
rect 81142 21734 81156 21786
rect 81180 21734 81194 21786
rect 81194 21734 81206 21786
rect 81206 21734 81236 21786
rect 81260 21734 81270 21786
rect 81270 21734 81316 21786
rect 81020 21732 81076 21734
rect 81100 21732 81156 21734
rect 81180 21732 81236 21734
rect 81260 21732 81316 21734
rect 62670 2352 62726 2408
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 65706 2352 65762 2408
rect 81020 20698 81076 20700
rect 81100 20698 81156 20700
rect 81180 20698 81236 20700
rect 81260 20698 81316 20700
rect 81020 20646 81066 20698
rect 81066 20646 81076 20698
rect 81100 20646 81130 20698
rect 81130 20646 81142 20698
rect 81142 20646 81156 20698
rect 81180 20646 81194 20698
rect 81194 20646 81206 20698
rect 81206 20646 81236 20698
rect 81260 20646 81270 20698
rect 81270 20646 81316 20698
rect 81020 20644 81076 20646
rect 81100 20644 81156 20646
rect 81180 20644 81236 20646
rect 81260 20644 81316 20646
rect 81020 19610 81076 19612
rect 81100 19610 81156 19612
rect 81180 19610 81236 19612
rect 81260 19610 81316 19612
rect 81020 19558 81066 19610
rect 81066 19558 81076 19610
rect 81100 19558 81130 19610
rect 81130 19558 81142 19610
rect 81142 19558 81156 19610
rect 81180 19558 81194 19610
rect 81194 19558 81206 19610
rect 81206 19558 81236 19610
rect 81260 19558 81270 19610
rect 81270 19558 81316 19610
rect 81020 19556 81076 19558
rect 81100 19556 81156 19558
rect 81180 19556 81236 19558
rect 81260 19556 81316 19558
rect 81020 18522 81076 18524
rect 81100 18522 81156 18524
rect 81180 18522 81236 18524
rect 81260 18522 81316 18524
rect 81020 18470 81066 18522
rect 81066 18470 81076 18522
rect 81100 18470 81130 18522
rect 81130 18470 81142 18522
rect 81142 18470 81156 18522
rect 81180 18470 81194 18522
rect 81194 18470 81206 18522
rect 81206 18470 81236 18522
rect 81260 18470 81270 18522
rect 81270 18470 81316 18522
rect 81020 18468 81076 18470
rect 81100 18468 81156 18470
rect 81180 18468 81236 18470
rect 81260 18468 81316 18470
rect 81020 17434 81076 17436
rect 81100 17434 81156 17436
rect 81180 17434 81236 17436
rect 81260 17434 81316 17436
rect 81020 17382 81066 17434
rect 81066 17382 81076 17434
rect 81100 17382 81130 17434
rect 81130 17382 81142 17434
rect 81142 17382 81156 17434
rect 81180 17382 81194 17434
rect 81194 17382 81206 17434
rect 81206 17382 81236 17434
rect 81260 17382 81270 17434
rect 81270 17382 81316 17434
rect 81020 17380 81076 17382
rect 81100 17380 81156 17382
rect 81180 17380 81236 17382
rect 81260 17380 81316 17382
rect 81020 16346 81076 16348
rect 81100 16346 81156 16348
rect 81180 16346 81236 16348
rect 81260 16346 81316 16348
rect 81020 16294 81066 16346
rect 81066 16294 81076 16346
rect 81100 16294 81130 16346
rect 81130 16294 81142 16346
rect 81142 16294 81156 16346
rect 81180 16294 81194 16346
rect 81194 16294 81206 16346
rect 81206 16294 81236 16346
rect 81260 16294 81270 16346
rect 81270 16294 81316 16346
rect 81020 16292 81076 16294
rect 81100 16292 81156 16294
rect 81180 16292 81236 16294
rect 81260 16292 81316 16294
rect 81020 15258 81076 15260
rect 81100 15258 81156 15260
rect 81180 15258 81236 15260
rect 81260 15258 81316 15260
rect 81020 15206 81066 15258
rect 81066 15206 81076 15258
rect 81100 15206 81130 15258
rect 81130 15206 81142 15258
rect 81142 15206 81156 15258
rect 81180 15206 81194 15258
rect 81194 15206 81206 15258
rect 81206 15206 81236 15258
rect 81260 15206 81270 15258
rect 81270 15206 81316 15258
rect 81020 15204 81076 15206
rect 81100 15204 81156 15206
rect 81180 15204 81236 15206
rect 81260 15204 81316 15206
rect 81020 14170 81076 14172
rect 81100 14170 81156 14172
rect 81180 14170 81236 14172
rect 81260 14170 81316 14172
rect 81020 14118 81066 14170
rect 81066 14118 81076 14170
rect 81100 14118 81130 14170
rect 81130 14118 81142 14170
rect 81142 14118 81156 14170
rect 81180 14118 81194 14170
rect 81194 14118 81206 14170
rect 81206 14118 81236 14170
rect 81260 14118 81270 14170
rect 81270 14118 81316 14170
rect 81020 14116 81076 14118
rect 81100 14116 81156 14118
rect 81180 14116 81236 14118
rect 81260 14116 81316 14118
rect 81020 13082 81076 13084
rect 81100 13082 81156 13084
rect 81180 13082 81236 13084
rect 81260 13082 81316 13084
rect 81020 13030 81066 13082
rect 81066 13030 81076 13082
rect 81100 13030 81130 13082
rect 81130 13030 81142 13082
rect 81142 13030 81156 13082
rect 81180 13030 81194 13082
rect 81194 13030 81206 13082
rect 81206 13030 81236 13082
rect 81260 13030 81270 13082
rect 81270 13030 81316 13082
rect 81020 13028 81076 13030
rect 81100 13028 81156 13030
rect 81180 13028 81236 13030
rect 81260 13028 81316 13030
rect 81020 11994 81076 11996
rect 81100 11994 81156 11996
rect 81180 11994 81236 11996
rect 81260 11994 81316 11996
rect 81020 11942 81066 11994
rect 81066 11942 81076 11994
rect 81100 11942 81130 11994
rect 81130 11942 81142 11994
rect 81142 11942 81156 11994
rect 81180 11942 81194 11994
rect 81194 11942 81206 11994
rect 81206 11942 81236 11994
rect 81260 11942 81270 11994
rect 81270 11942 81316 11994
rect 81020 11940 81076 11942
rect 81100 11940 81156 11942
rect 81180 11940 81236 11942
rect 81260 11940 81316 11942
rect 81020 10906 81076 10908
rect 81100 10906 81156 10908
rect 81180 10906 81236 10908
rect 81260 10906 81316 10908
rect 81020 10854 81066 10906
rect 81066 10854 81076 10906
rect 81100 10854 81130 10906
rect 81130 10854 81142 10906
rect 81142 10854 81156 10906
rect 81180 10854 81194 10906
rect 81194 10854 81206 10906
rect 81206 10854 81236 10906
rect 81260 10854 81270 10906
rect 81270 10854 81316 10906
rect 81020 10852 81076 10854
rect 81100 10852 81156 10854
rect 81180 10852 81236 10854
rect 81260 10852 81316 10854
rect 81020 9818 81076 9820
rect 81100 9818 81156 9820
rect 81180 9818 81236 9820
rect 81260 9818 81316 9820
rect 81020 9766 81066 9818
rect 81066 9766 81076 9818
rect 81100 9766 81130 9818
rect 81130 9766 81142 9818
rect 81142 9766 81156 9818
rect 81180 9766 81194 9818
rect 81194 9766 81206 9818
rect 81206 9766 81236 9818
rect 81260 9766 81270 9818
rect 81270 9766 81316 9818
rect 81020 9764 81076 9766
rect 81100 9764 81156 9766
rect 81180 9764 81236 9766
rect 81260 9764 81316 9766
rect 81020 8730 81076 8732
rect 81100 8730 81156 8732
rect 81180 8730 81236 8732
rect 81260 8730 81316 8732
rect 81020 8678 81066 8730
rect 81066 8678 81076 8730
rect 81100 8678 81130 8730
rect 81130 8678 81142 8730
rect 81142 8678 81156 8730
rect 81180 8678 81194 8730
rect 81194 8678 81206 8730
rect 81206 8678 81236 8730
rect 81260 8678 81270 8730
rect 81270 8678 81316 8730
rect 81020 8676 81076 8678
rect 81100 8676 81156 8678
rect 81180 8676 81236 8678
rect 81260 8676 81316 8678
rect 81020 7642 81076 7644
rect 81100 7642 81156 7644
rect 81180 7642 81236 7644
rect 81260 7642 81316 7644
rect 81020 7590 81066 7642
rect 81066 7590 81076 7642
rect 81100 7590 81130 7642
rect 81130 7590 81142 7642
rect 81142 7590 81156 7642
rect 81180 7590 81194 7642
rect 81194 7590 81206 7642
rect 81206 7590 81236 7642
rect 81260 7590 81270 7642
rect 81270 7590 81316 7642
rect 81020 7588 81076 7590
rect 81100 7588 81156 7590
rect 81180 7588 81236 7590
rect 81260 7588 81316 7590
rect 81020 6554 81076 6556
rect 81100 6554 81156 6556
rect 81180 6554 81236 6556
rect 81260 6554 81316 6556
rect 81020 6502 81066 6554
rect 81066 6502 81076 6554
rect 81100 6502 81130 6554
rect 81130 6502 81142 6554
rect 81142 6502 81156 6554
rect 81180 6502 81194 6554
rect 81194 6502 81206 6554
rect 81206 6502 81236 6554
rect 81260 6502 81270 6554
rect 81270 6502 81316 6554
rect 81020 6500 81076 6502
rect 81100 6500 81156 6502
rect 81180 6500 81236 6502
rect 81260 6500 81316 6502
rect 81020 5466 81076 5468
rect 81100 5466 81156 5468
rect 81180 5466 81236 5468
rect 81260 5466 81316 5468
rect 81020 5414 81066 5466
rect 81066 5414 81076 5466
rect 81100 5414 81130 5466
rect 81130 5414 81142 5466
rect 81142 5414 81156 5466
rect 81180 5414 81194 5466
rect 81194 5414 81206 5466
rect 81206 5414 81236 5466
rect 81260 5414 81270 5466
rect 81270 5414 81316 5466
rect 81020 5412 81076 5414
rect 81100 5412 81156 5414
rect 81180 5412 81236 5414
rect 81260 5412 81316 5414
rect 81020 4378 81076 4380
rect 81100 4378 81156 4380
rect 81180 4378 81236 4380
rect 81260 4378 81316 4380
rect 81020 4326 81066 4378
rect 81066 4326 81076 4378
rect 81100 4326 81130 4378
rect 81130 4326 81142 4378
rect 81142 4326 81156 4378
rect 81180 4326 81194 4378
rect 81194 4326 81206 4378
rect 81206 4326 81236 4378
rect 81260 4326 81270 4378
rect 81270 4326 81316 4378
rect 81020 4324 81076 4326
rect 81100 4324 81156 4326
rect 81180 4324 81236 4326
rect 81260 4324 81316 4326
rect 81020 3290 81076 3292
rect 81100 3290 81156 3292
rect 81180 3290 81236 3292
rect 81260 3290 81316 3292
rect 81020 3238 81066 3290
rect 81066 3238 81076 3290
rect 81100 3238 81130 3290
rect 81130 3238 81142 3290
rect 81142 3238 81156 3290
rect 81180 3238 81194 3290
rect 81194 3238 81206 3290
rect 81206 3238 81236 3290
rect 81260 3238 81270 3290
rect 81270 3238 81316 3290
rect 81020 3236 81076 3238
rect 81100 3236 81156 3238
rect 81180 3236 81236 3238
rect 81260 3236 81316 3238
rect 81020 2202 81076 2204
rect 81100 2202 81156 2204
rect 81180 2202 81236 2204
rect 81260 2202 81316 2204
rect 81020 2150 81066 2202
rect 81066 2150 81076 2202
rect 81100 2150 81130 2202
rect 81130 2150 81142 2202
rect 81142 2150 81156 2202
rect 81180 2150 81194 2202
rect 81194 2150 81206 2202
rect 81206 2150 81236 2202
rect 81260 2150 81270 2202
rect 81270 2150 81316 2202
rect 81020 2148 81076 2150
rect 81100 2148 81156 2150
rect 81180 2148 81236 2150
rect 81260 2148 81316 2150
rect 96380 37562 96436 37564
rect 96460 37562 96516 37564
rect 96540 37562 96596 37564
rect 96620 37562 96676 37564
rect 96380 37510 96426 37562
rect 96426 37510 96436 37562
rect 96460 37510 96490 37562
rect 96490 37510 96502 37562
rect 96502 37510 96516 37562
rect 96540 37510 96554 37562
rect 96554 37510 96566 37562
rect 96566 37510 96596 37562
rect 96620 37510 96630 37562
rect 96630 37510 96676 37562
rect 96380 37508 96436 37510
rect 96460 37508 96516 37510
rect 96540 37508 96596 37510
rect 96620 37508 96676 37510
rect 96380 36474 96436 36476
rect 96460 36474 96516 36476
rect 96540 36474 96596 36476
rect 96620 36474 96676 36476
rect 96380 36422 96426 36474
rect 96426 36422 96436 36474
rect 96460 36422 96490 36474
rect 96490 36422 96502 36474
rect 96502 36422 96516 36474
rect 96540 36422 96554 36474
rect 96554 36422 96566 36474
rect 96566 36422 96596 36474
rect 96620 36422 96630 36474
rect 96630 36422 96676 36474
rect 96380 36420 96436 36422
rect 96460 36420 96516 36422
rect 96540 36420 96596 36422
rect 96620 36420 96676 36422
rect 96380 35386 96436 35388
rect 96460 35386 96516 35388
rect 96540 35386 96596 35388
rect 96620 35386 96676 35388
rect 96380 35334 96426 35386
rect 96426 35334 96436 35386
rect 96460 35334 96490 35386
rect 96490 35334 96502 35386
rect 96502 35334 96516 35386
rect 96540 35334 96554 35386
rect 96554 35334 96566 35386
rect 96566 35334 96596 35386
rect 96620 35334 96630 35386
rect 96630 35334 96676 35386
rect 96380 35332 96436 35334
rect 96460 35332 96516 35334
rect 96540 35332 96596 35334
rect 96620 35332 96676 35334
rect 96380 34298 96436 34300
rect 96460 34298 96516 34300
rect 96540 34298 96596 34300
rect 96620 34298 96676 34300
rect 96380 34246 96426 34298
rect 96426 34246 96436 34298
rect 96460 34246 96490 34298
rect 96490 34246 96502 34298
rect 96502 34246 96516 34298
rect 96540 34246 96554 34298
rect 96554 34246 96566 34298
rect 96566 34246 96596 34298
rect 96620 34246 96630 34298
rect 96630 34246 96676 34298
rect 96380 34244 96436 34246
rect 96460 34244 96516 34246
rect 96540 34244 96596 34246
rect 96620 34244 96676 34246
rect 96380 33210 96436 33212
rect 96460 33210 96516 33212
rect 96540 33210 96596 33212
rect 96620 33210 96676 33212
rect 96380 33158 96426 33210
rect 96426 33158 96436 33210
rect 96460 33158 96490 33210
rect 96490 33158 96502 33210
rect 96502 33158 96516 33210
rect 96540 33158 96554 33210
rect 96554 33158 96566 33210
rect 96566 33158 96596 33210
rect 96620 33158 96630 33210
rect 96630 33158 96676 33210
rect 96380 33156 96436 33158
rect 96460 33156 96516 33158
rect 96540 33156 96596 33158
rect 96620 33156 96676 33158
rect 96380 32122 96436 32124
rect 96460 32122 96516 32124
rect 96540 32122 96596 32124
rect 96620 32122 96676 32124
rect 96380 32070 96426 32122
rect 96426 32070 96436 32122
rect 96460 32070 96490 32122
rect 96490 32070 96502 32122
rect 96502 32070 96516 32122
rect 96540 32070 96554 32122
rect 96554 32070 96566 32122
rect 96566 32070 96596 32122
rect 96620 32070 96630 32122
rect 96630 32070 96676 32122
rect 96380 32068 96436 32070
rect 96460 32068 96516 32070
rect 96540 32068 96596 32070
rect 96620 32068 96676 32070
rect 96380 31034 96436 31036
rect 96460 31034 96516 31036
rect 96540 31034 96596 31036
rect 96620 31034 96676 31036
rect 96380 30982 96426 31034
rect 96426 30982 96436 31034
rect 96460 30982 96490 31034
rect 96490 30982 96502 31034
rect 96502 30982 96516 31034
rect 96540 30982 96554 31034
rect 96554 30982 96566 31034
rect 96566 30982 96596 31034
rect 96620 30982 96630 31034
rect 96630 30982 96676 31034
rect 96380 30980 96436 30982
rect 96460 30980 96516 30982
rect 96540 30980 96596 30982
rect 96620 30980 96676 30982
rect 96380 29946 96436 29948
rect 96460 29946 96516 29948
rect 96540 29946 96596 29948
rect 96620 29946 96676 29948
rect 96380 29894 96426 29946
rect 96426 29894 96436 29946
rect 96460 29894 96490 29946
rect 96490 29894 96502 29946
rect 96502 29894 96516 29946
rect 96540 29894 96554 29946
rect 96554 29894 96566 29946
rect 96566 29894 96596 29946
rect 96620 29894 96630 29946
rect 96630 29894 96676 29946
rect 96380 29892 96436 29894
rect 96460 29892 96516 29894
rect 96540 29892 96596 29894
rect 96620 29892 96676 29894
rect 96380 28858 96436 28860
rect 96460 28858 96516 28860
rect 96540 28858 96596 28860
rect 96620 28858 96676 28860
rect 96380 28806 96426 28858
rect 96426 28806 96436 28858
rect 96460 28806 96490 28858
rect 96490 28806 96502 28858
rect 96502 28806 96516 28858
rect 96540 28806 96554 28858
rect 96554 28806 96566 28858
rect 96566 28806 96596 28858
rect 96620 28806 96630 28858
rect 96630 28806 96676 28858
rect 96380 28804 96436 28806
rect 96460 28804 96516 28806
rect 96540 28804 96596 28806
rect 96620 28804 96676 28806
rect 96380 27770 96436 27772
rect 96460 27770 96516 27772
rect 96540 27770 96596 27772
rect 96620 27770 96676 27772
rect 96380 27718 96426 27770
rect 96426 27718 96436 27770
rect 96460 27718 96490 27770
rect 96490 27718 96502 27770
rect 96502 27718 96516 27770
rect 96540 27718 96554 27770
rect 96554 27718 96566 27770
rect 96566 27718 96596 27770
rect 96620 27718 96630 27770
rect 96630 27718 96676 27770
rect 96380 27716 96436 27718
rect 96460 27716 96516 27718
rect 96540 27716 96596 27718
rect 96620 27716 96676 27718
rect 96380 26682 96436 26684
rect 96460 26682 96516 26684
rect 96540 26682 96596 26684
rect 96620 26682 96676 26684
rect 96380 26630 96426 26682
rect 96426 26630 96436 26682
rect 96460 26630 96490 26682
rect 96490 26630 96502 26682
rect 96502 26630 96516 26682
rect 96540 26630 96554 26682
rect 96554 26630 96566 26682
rect 96566 26630 96596 26682
rect 96620 26630 96630 26682
rect 96630 26630 96676 26682
rect 96380 26628 96436 26630
rect 96460 26628 96516 26630
rect 96540 26628 96596 26630
rect 96620 26628 96676 26630
rect 96380 25594 96436 25596
rect 96460 25594 96516 25596
rect 96540 25594 96596 25596
rect 96620 25594 96676 25596
rect 96380 25542 96426 25594
rect 96426 25542 96436 25594
rect 96460 25542 96490 25594
rect 96490 25542 96502 25594
rect 96502 25542 96516 25594
rect 96540 25542 96554 25594
rect 96554 25542 96566 25594
rect 96566 25542 96596 25594
rect 96620 25542 96630 25594
rect 96630 25542 96676 25594
rect 96380 25540 96436 25542
rect 96460 25540 96516 25542
rect 96540 25540 96596 25542
rect 96620 25540 96676 25542
rect 96380 24506 96436 24508
rect 96460 24506 96516 24508
rect 96540 24506 96596 24508
rect 96620 24506 96676 24508
rect 96380 24454 96426 24506
rect 96426 24454 96436 24506
rect 96460 24454 96490 24506
rect 96490 24454 96502 24506
rect 96502 24454 96516 24506
rect 96540 24454 96554 24506
rect 96554 24454 96566 24506
rect 96566 24454 96596 24506
rect 96620 24454 96630 24506
rect 96630 24454 96676 24506
rect 96380 24452 96436 24454
rect 96460 24452 96516 24454
rect 96540 24452 96596 24454
rect 96620 24452 96676 24454
rect 96380 23418 96436 23420
rect 96460 23418 96516 23420
rect 96540 23418 96596 23420
rect 96620 23418 96676 23420
rect 96380 23366 96426 23418
rect 96426 23366 96436 23418
rect 96460 23366 96490 23418
rect 96490 23366 96502 23418
rect 96502 23366 96516 23418
rect 96540 23366 96554 23418
rect 96554 23366 96566 23418
rect 96566 23366 96596 23418
rect 96620 23366 96630 23418
rect 96630 23366 96676 23418
rect 96380 23364 96436 23366
rect 96460 23364 96516 23366
rect 96540 23364 96596 23366
rect 96620 23364 96676 23366
rect 96380 22330 96436 22332
rect 96460 22330 96516 22332
rect 96540 22330 96596 22332
rect 96620 22330 96676 22332
rect 96380 22278 96426 22330
rect 96426 22278 96436 22330
rect 96460 22278 96490 22330
rect 96490 22278 96502 22330
rect 96502 22278 96516 22330
rect 96540 22278 96554 22330
rect 96554 22278 96566 22330
rect 96566 22278 96596 22330
rect 96620 22278 96630 22330
rect 96630 22278 96676 22330
rect 96380 22276 96436 22278
rect 96460 22276 96516 22278
rect 96540 22276 96596 22278
rect 96620 22276 96676 22278
rect 96380 21242 96436 21244
rect 96460 21242 96516 21244
rect 96540 21242 96596 21244
rect 96620 21242 96676 21244
rect 96380 21190 96426 21242
rect 96426 21190 96436 21242
rect 96460 21190 96490 21242
rect 96490 21190 96502 21242
rect 96502 21190 96516 21242
rect 96540 21190 96554 21242
rect 96554 21190 96566 21242
rect 96566 21190 96596 21242
rect 96620 21190 96630 21242
rect 96630 21190 96676 21242
rect 96380 21188 96436 21190
rect 96460 21188 96516 21190
rect 96540 21188 96596 21190
rect 96620 21188 96676 21190
rect 96380 20154 96436 20156
rect 96460 20154 96516 20156
rect 96540 20154 96596 20156
rect 96620 20154 96676 20156
rect 96380 20102 96426 20154
rect 96426 20102 96436 20154
rect 96460 20102 96490 20154
rect 96490 20102 96502 20154
rect 96502 20102 96516 20154
rect 96540 20102 96554 20154
rect 96554 20102 96566 20154
rect 96566 20102 96596 20154
rect 96620 20102 96630 20154
rect 96630 20102 96676 20154
rect 96380 20100 96436 20102
rect 96460 20100 96516 20102
rect 96540 20100 96596 20102
rect 96620 20100 96676 20102
rect 96380 19066 96436 19068
rect 96460 19066 96516 19068
rect 96540 19066 96596 19068
rect 96620 19066 96676 19068
rect 96380 19014 96426 19066
rect 96426 19014 96436 19066
rect 96460 19014 96490 19066
rect 96490 19014 96502 19066
rect 96502 19014 96516 19066
rect 96540 19014 96554 19066
rect 96554 19014 96566 19066
rect 96566 19014 96596 19066
rect 96620 19014 96630 19066
rect 96630 19014 96676 19066
rect 96380 19012 96436 19014
rect 96460 19012 96516 19014
rect 96540 19012 96596 19014
rect 96620 19012 96676 19014
rect 96380 17978 96436 17980
rect 96460 17978 96516 17980
rect 96540 17978 96596 17980
rect 96620 17978 96676 17980
rect 96380 17926 96426 17978
rect 96426 17926 96436 17978
rect 96460 17926 96490 17978
rect 96490 17926 96502 17978
rect 96502 17926 96516 17978
rect 96540 17926 96554 17978
rect 96554 17926 96566 17978
rect 96566 17926 96596 17978
rect 96620 17926 96630 17978
rect 96630 17926 96676 17978
rect 96380 17924 96436 17926
rect 96460 17924 96516 17926
rect 96540 17924 96596 17926
rect 96620 17924 96676 17926
rect 96380 16890 96436 16892
rect 96460 16890 96516 16892
rect 96540 16890 96596 16892
rect 96620 16890 96676 16892
rect 96380 16838 96426 16890
rect 96426 16838 96436 16890
rect 96460 16838 96490 16890
rect 96490 16838 96502 16890
rect 96502 16838 96516 16890
rect 96540 16838 96554 16890
rect 96554 16838 96566 16890
rect 96566 16838 96596 16890
rect 96620 16838 96630 16890
rect 96630 16838 96676 16890
rect 96380 16836 96436 16838
rect 96460 16836 96516 16838
rect 96540 16836 96596 16838
rect 96620 16836 96676 16838
rect 96380 15802 96436 15804
rect 96460 15802 96516 15804
rect 96540 15802 96596 15804
rect 96620 15802 96676 15804
rect 96380 15750 96426 15802
rect 96426 15750 96436 15802
rect 96460 15750 96490 15802
rect 96490 15750 96502 15802
rect 96502 15750 96516 15802
rect 96540 15750 96554 15802
rect 96554 15750 96566 15802
rect 96566 15750 96596 15802
rect 96620 15750 96630 15802
rect 96630 15750 96676 15802
rect 96380 15748 96436 15750
rect 96460 15748 96516 15750
rect 96540 15748 96596 15750
rect 96620 15748 96676 15750
rect 96380 14714 96436 14716
rect 96460 14714 96516 14716
rect 96540 14714 96596 14716
rect 96620 14714 96676 14716
rect 96380 14662 96426 14714
rect 96426 14662 96436 14714
rect 96460 14662 96490 14714
rect 96490 14662 96502 14714
rect 96502 14662 96516 14714
rect 96540 14662 96554 14714
rect 96554 14662 96566 14714
rect 96566 14662 96596 14714
rect 96620 14662 96630 14714
rect 96630 14662 96676 14714
rect 96380 14660 96436 14662
rect 96460 14660 96516 14662
rect 96540 14660 96596 14662
rect 96620 14660 96676 14662
rect 96380 13626 96436 13628
rect 96460 13626 96516 13628
rect 96540 13626 96596 13628
rect 96620 13626 96676 13628
rect 96380 13574 96426 13626
rect 96426 13574 96436 13626
rect 96460 13574 96490 13626
rect 96490 13574 96502 13626
rect 96502 13574 96516 13626
rect 96540 13574 96554 13626
rect 96554 13574 96566 13626
rect 96566 13574 96596 13626
rect 96620 13574 96630 13626
rect 96630 13574 96676 13626
rect 96380 13572 96436 13574
rect 96460 13572 96516 13574
rect 96540 13572 96596 13574
rect 96620 13572 96676 13574
rect 96380 12538 96436 12540
rect 96460 12538 96516 12540
rect 96540 12538 96596 12540
rect 96620 12538 96676 12540
rect 96380 12486 96426 12538
rect 96426 12486 96436 12538
rect 96460 12486 96490 12538
rect 96490 12486 96502 12538
rect 96502 12486 96516 12538
rect 96540 12486 96554 12538
rect 96554 12486 96566 12538
rect 96566 12486 96596 12538
rect 96620 12486 96630 12538
rect 96630 12486 96676 12538
rect 96380 12484 96436 12486
rect 96460 12484 96516 12486
rect 96540 12484 96596 12486
rect 96620 12484 96676 12486
rect 96380 11450 96436 11452
rect 96460 11450 96516 11452
rect 96540 11450 96596 11452
rect 96620 11450 96676 11452
rect 96380 11398 96426 11450
rect 96426 11398 96436 11450
rect 96460 11398 96490 11450
rect 96490 11398 96502 11450
rect 96502 11398 96516 11450
rect 96540 11398 96554 11450
rect 96554 11398 96566 11450
rect 96566 11398 96596 11450
rect 96620 11398 96630 11450
rect 96630 11398 96676 11450
rect 96380 11396 96436 11398
rect 96460 11396 96516 11398
rect 96540 11396 96596 11398
rect 96620 11396 96676 11398
rect 96380 10362 96436 10364
rect 96460 10362 96516 10364
rect 96540 10362 96596 10364
rect 96620 10362 96676 10364
rect 96380 10310 96426 10362
rect 96426 10310 96436 10362
rect 96460 10310 96490 10362
rect 96490 10310 96502 10362
rect 96502 10310 96516 10362
rect 96540 10310 96554 10362
rect 96554 10310 96566 10362
rect 96566 10310 96596 10362
rect 96620 10310 96630 10362
rect 96630 10310 96676 10362
rect 96380 10308 96436 10310
rect 96460 10308 96516 10310
rect 96540 10308 96596 10310
rect 96620 10308 96676 10310
rect 96380 9274 96436 9276
rect 96460 9274 96516 9276
rect 96540 9274 96596 9276
rect 96620 9274 96676 9276
rect 96380 9222 96426 9274
rect 96426 9222 96436 9274
rect 96460 9222 96490 9274
rect 96490 9222 96502 9274
rect 96502 9222 96516 9274
rect 96540 9222 96554 9274
rect 96554 9222 96566 9274
rect 96566 9222 96596 9274
rect 96620 9222 96630 9274
rect 96630 9222 96676 9274
rect 96380 9220 96436 9222
rect 96460 9220 96516 9222
rect 96540 9220 96596 9222
rect 96620 9220 96676 9222
rect 96380 8186 96436 8188
rect 96460 8186 96516 8188
rect 96540 8186 96596 8188
rect 96620 8186 96676 8188
rect 96380 8134 96426 8186
rect 96426 8134 96436 8186
rect 96460 8134 96490 8186
rect 96490 8134 96502 8186
rect 96502 8134 96516 8186
rect 96540 8134 96554 8186
rect 96554 8134 96566 8186
rect 96566 8134 96596 8186
rect 96620 8134 96630 8186
rect 96630 8134 96676 8186
rect 96380 8132 96436 8134
rect 96460 8132 96516 8134
rect 96540 8132 96596 8134
rect 96620 8132 96676 8134
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 104254 2896 104310 2952
rect 111740 37018 111796 37020
rect 111820 37018 111876 37020
rect 111900 37018 111956 37020
rect 111980 37018 112036 37020
rect 111740 36966 111786 37018
rect 111786 36966 111796 37018
rect 111820 36966 111850 37018
rect 111850 36966 111862 37018
rect 111862 36966 111876 37018
rect 111900 36966 111914 37018
rect 111914 36966 111926 37018
rect 111926 36966 111956 37018
rect 111980 36966 111990 37018
rect 111990 36966 112036 37018
rect 111740 36964 111796 36966
rect 111820 36964 111876 36966
rect 111900 36964 111956 36966
rect 111980 36964 112036 36966
rect 111740 35930 111796 35932
rect 111820 35930 111876 35932
rect 111900 35930 111956 35932
rect 111980 35930 112036 35932
rect 111740 35878 111786 35930
rect 111786 35878 111796 35930
rect 111820 35878 111850 35930
rect 111850 35878 111862 35930
rect 111862 35878 111876 35930
rect 111900 35878 111914 35930
rect 111914 35878 111926 35930
rect 111926 35878 111956 35930
rect 111980 35878 111990 35930
rect 111990 35878 112036 35930
rect 111740 35876 111796 35878
rect 111820 35876 111876 35878
rect 111900 35876 111956 35878
rect 111980 35876 112036 35878
rect 111740 34842 111796 34844
rect 111820 34842 111876 34844
rect 111900 34842 111956 34844
rect 111980 34842 112036 34844
rect 111740 34790 111786 34842
rect 111786 34790 111796 34842
rect 111820 34790 111850 34842
rect 111850 34790 111862 34842
rect 111862 34790 111876 34842
rect 111900 34790 111914 34842
rect 111914 34790 111926 34842
rect 111926 34790 111956 34842
rect 111980 34790 111990 34842
rect 111990 34790 112036 34842
rect 111740 34788 111796 34790
rect 111820 34788 111876 34790
rect 111900 34788 111956 34790
rect 111980 34788 112036 34790
rect 111740 33754 111796 33756
rect 111820 33754 111876 33756
rect 111900 33754 111956 33756
rect 111980 33754 112036 33756
rect 111740 33702 111786 33754
rect 111786 33702 111796 33754
rect 111820 33702 111850 33754
rect 111850 33702 111862 33754
rect 111862 33702 111876 33754
rect 111900 33702 111914 33754
rect 111914 33702 111926 33754
rect 111926 33702 111956 33754
rect 111980 33702 111990 33754
rect 111990 33702 112036 33754
rect 111740 33700 111796 33702
rect 111820 33700 111876 33702
rect 111900 33700 111956 33702
rect 111980 33700 112036 33702
rect 111740 32666 111796 32668
rect 111820 32666 111876 32668
rect 111900 32666 111956 32668
rect 111980 32666 112036 32668
rect 111740 32614 111786 32666
rect 111786 32614 111796 32666
rect 111820 32614 111850 32666
rect 111850 32614 111862 32666
rect 111862 32614 111876 32666
rect 111900 32614 111914 32666
rect 111914 32614 111926 32666
rect 111926 32614 111956 32666
rect 111980 32614 111990 32666
rect 111990 32614 112036 32666
rect 111740 32612 111796 32614
rect 111820 32612 111876 32614
rect 111900 32612 111956 32614
rect 111980 32612 112036 32614
rect 111740 31578 111796 31580
rect 111820 31578 111876 31580
rect 111900 31578 111956 31580
rect 111980 31578 112036 31580
rect 111740 31526 111786 31578
rect 111786 31526 111796 31578
rect 111820 31526 111850 31578
rect 111850 31526 111862 31578
rect 111862 31526 111876 31578
rect 111900 31526 111914 31578
rect 111914 31526 111926 31578
rect 111926 31526 111956 31578
rect 111980 31526 111990 31578
rect 111990 31526 112036 31578
rect 111740 31524 111796 31526
rect 111820 31524 111876 31526
rect 111900 31524 111956 31526
rect 111980 31524 112036 31526
rect 111740 30490 111796 30492
rect 111820 30490 111876 30492
rect 111900 30490 111956 30492
rect 111980 30490 112036 30492
rect 111740 30438 111786 30490
rect 111786 30438 111796 30490
rect 111820 30438 111850 30490
rect 111850 30438 111862 30490
rect 111862 30438 111876 30490
rect 111900 30438 111914 30490
rect 111914 30438 111926 30490
rect 111926 30438 111956 30490
rect 111980 30438 111990 30490
rect 111990 30438 112036 30490
rect 111740 30436 111796 30438
rect 111820 30436 111876 30438
rect 111900 30436 111956 30438
rect 111980 30436 112036 30438
rect 111740 29402 111796 29404
rect 111820 29402 111876 29404
rect 111900 29402 111956 29404
rect 111980 29402 112036 29404
rect 111740 29350 111786 29402
rect 111786 29350 111796 29402
rect 111820 29350 111850 29402
rect 111850 29350 111862 29402
rect 111862 29350 111876 29402
rect 111900 29350 111914 29402
rect 111914 29350 111926 29402
rect 111926 29350 111956 29402
rect 111980 29350 111990 29402
rect 111990 29350 112036 29402
rect 111740 29348 111796 29350
rect 111820 29348 111876 29350
rect 111900 29348 111956 29350
rect 111980 29348 112036 29350
rect 111740 28314 111796 28316
rect 111820 28314 111876 28316
rect 111900 28314 111956 28316
rect 111980 28314 112036 28316
rect 111740 28262 111786 28314
rect 111786 28262 111796 28314
rect 111820 28262 111850 28314
rect 111850 28262 111862 28314
rect 111862 28262 111876 28314
rect 111900 28262 111914 28314
rect 111914 28262 111926 28314
rect 111926 28262 111956 28314
rect 111980 28262 111990 28314
rect 111990 28262 112036 28314
rect 111740 28260 111796 28262
rect 111820 28260 111876 28262
rect 111900 28260 111956 28262
rect 111980 28260 112036 28262
rect 111740 27226 111796 27228
rect 111820 27226 111876 27228
rect 111900 27226 111956 27228
rect 111980 27226 112036 27228
rect 111740 27174 111786 27226
rect 111786 27174 111796 27226
rect 111820 27174 111850 27226
rect 111850 27174 111862 27226
rect 111862 27174 111876 27226
rect 111900 27174 111914 27226
rect 111914 27174 111926 27226
rect 111926 27174 111956 27226
rect 111980 27174 111990 27226
rect 111990 27174 112036 27226
rect 111740 27172 111796 27174
rect 111820 27172 111876 27174
rect 111900 27172 111956 27174
rect 111980 27172 112036 27174
rect 111740 26138 111796 26140
rect 111820 26138 111876 26140
rect 111900 26138 111956 26140
rect 111980 26138 112036 26140
rect 111740 26086 111786 26138
rect 111786 26086 111796 26138
rect 111820 26086 111850 26138
rect 111850 26086 111862 26138
rect 111862 26086 111876 26138
rect 111900 26086 111914 26138
rect 111914 26086 111926 26138
rect 111926 26086 111956 26138
rect 111980 26086 111990 26138
rect 111990 26086 112036 26138
rect 111740 26084 111796 26086
rect 111820 26084 111876 26086
rect 111900 26084 111956 26086
rect 111980 26084 112036 26086
rect 111740 25050 111796 25052
rect 111820 25050 111876 25052
rect 111900 25050 111956 25052
rect 111980 25050 112036 25052
rect 111740 24998 111786 25050
rect 111786 24998 111796 25050
rect 111820 24998 111850 25050
rect 111850 24998 111862 25050
rect 111862 24998 111876 25050
rect 111900 24998 111914 25050
rect 111914 24998 111926 25050
rect 111926 24998 111956 25050
rect 111980 24998 111990 25050
rect 111990 24998 112036 25050
rect 111740 24996 111796 24998
rect 111820 24996 111876 24998
rect 111900 24996 111956 24998
rect 111980 24996 112036 24998
rect 111740 23962 111796 23964
rect 111820 23962 111876 23964
rect 111900 23962 111956 23964
rect 111980 23962 112036 23964
rect 111740 23910 111786 23962
rect 111786 23910 111796 23962
rect 111820 23910 111850 23962
rect 111850 23910 111862 23962
rect 111862 23910 111876 23962
rect 111900 23910 111914 23962
rect 111914 23910 111926 23962
rect 111926 23910 111956 23962
rect 111980 23910 111990 23962
rect 111990 23910 112036 23962
rect 111740 23908 111796 23910
rect 111820 23908 111876 23910
rect 111900 23908 111956 23910
rect 111980 23908 112036 23910
rect 111740 22874 111796 22876
rect 111820 22874 111876 22876
rect 111900 22874 111956 22876
rect 111980 22874 112036 22876
rect 111740 22822 111786 22874
rect 111786 22822 111796 22874
rect 111820 22822 111850 22874
rect 111850 22822 111862 22874
rect 111862 22822 111876 22874
rect 111900 22822 111914 22874
rect 111914 22822 111926 22874
rect 111926 22822 111956 22874
rect 111980 22822 111990 22874
rect 111990 22822 112036 22874
rect 111740 22820 111796 22822
rect 111820 22820 111876 22822
rect 111900 22820 111956 22822
rect 111980 22820 112036 22822
rect 111740 21786 111796 21788
rect 111820 21786 111876 21788
rect 111900 21786 111956 21788
rect 111980 21786 112036 21788
rect 111740 21734 111786 21786
rect 111786 21734 111796 21786
rect 111820 21734 111850 21786
rect 111850 21734 111862 21786
rect 111862 21734 111876 21786
rect 111900 21734 111914 21786
rect 111914 21734 111926 21786
rect 111926 21734 111956 21786
rect 111980 21734 111990 21786
rect 111990 21734 112036 21786
rect 111740 21732 111796 21734
rect 111820 21732 111876 21734
rect 111900 21732 111956 21734
rect 111980 21732 112036 21734
rect 111740 20698 111796 20700
rect 111820 20698 111876 20700
rect 111900 20698 111956 20700
rect 111980 20698 112036 20700
rect 111740 20646 111786 20698
rect 111786 20646 111796 20698
rect 111820 20646 111850 20698
rect 111850 20646 111862 20698
rect 111862 20646 111876 20698
rect 111900 20646 111914 20698
rect 111914 20646 111926 20698
rect 111926 20646 111956 20698
rect 111980 20646 111990 20698
rect 111990 20646 112036 20698
rect 111740 20644 111796 20646
rect 111820 20644 111876 20646
rect 111900 20644 111956 20646
rect 111980 20644 112036 20646
rect 111740 19610 111796 19612
rect 111820 19610 111876 19612
rect 111900 19610 111956 19612
rect 111980 19610 112036 19612
rect 111740 19558 111786 19610
rect 111786 19558 111796 19610
rect 111820 19558 111850 19610
rect 111850 19558 111862 19610
rect 111862 19558 111876 19610
rect 111900 19558 111914 19610
rect 111914 19558 111926 19610
rect 111926 19558 111956 19610
rect 111980 19558 111990 19610
rect 111990 19558 112036 19610
rect 111740 19556 111796 19558
rect 111820 19556 111876 19558
rect 111900 19556 111956 19558
rect 111980 19556 112036 19558
rect 111740 18522 111796 18524
rect 111820 18522 111876 18524
rect 111900 18522 111956 18524
rect 111980 18522 112036 18524
rect 111740 18470 111786 18522
rect 111786 18470 111796 18522
rect 111820 18470 111850 18522
rect 111850 18470 111862 18522
rect 111862 18470 111876 18522
rect 111900 18470 111914 18522
rect 111914 18470 111926 18522
rect 111926 18470 111956 18522
rect 111980 18470 111990 18522
rect 111990 18470 112036 18522
rect 111740 18468 111796 18470
rect 111820 18468 111876 18470
rect 111900 18468 111956 18470
rect 111980 18468 112036 18470
rect 111740 17434 111796 17436
rect 111820 17434 111876 17436
rect 111900 17434 111956 17436
rect 111980 17434 112036 17436
rect 111740 17382 111786 17434
rect 111786 17382 111796 17434
rect 111820 17382 111850 17434
rect 111850 17382 111862 17434
rect 111862 17382 111876 17434
rect 111900 17382 111914 17434
rect 111914 17382 111926 17434
rect 111926 17382 111956 17434
rect 111980 17382 111990 17434
rect 111990 17382 112036 17434
rect 111740 17380 111796 17382
rect 111820 17380 111876 17382
rect 111900 17380 111956 17382
rect 111980 17380 112036 17382
rect 111740 16346 111796 16348
rect 111820 16346 111876 16348
rect 111900 16346 111956 16348
rect 111980 16346 112036 16348
rect 111740 16294 111786 16346
rect 111786 16294 111796 16346
rect 111820 16294 111850 16346
rect 111850 16294 111862 16346
rect 111862 16294 111876 16346
rect 111900 16294 111914 16346
rect 111914 16294 111926 16346
rect 111926 16294 111956 16346
rect 111980 16294 111990 16346
rect 111990 16294 112036 16346
rect 111740 16292 111796 16294
rect 111820 16292 111876 16294
rect 111900 16292 111956 16294
rect 111980 16292 112036 16294
rect 111740 15258 111796 15260
rect 111820 15258 111876 15260
rect 111900 15258 111956 15260
rect 111980 15258 112036 15260
rect 111740 15206 111786 15258
rect 111786 15206 111796 15258
rect 111820 15206 111850 15258
rect 111850 15206 111862 15258
rect 111862 15206 111876 15258
rect 111900 15206 111914 15258
rect 111914 15206 111926 15258
rect 111926 15206 111956 15258
rect 111980 15206 111990 15258
rect 111990 15206 112036 15258
rect 111740 15204 111796 15206
rect 111820 15204 111876 15206
rect 111900 15204 111956 15206
rect 111980 15204 112036 15206
rect 111740 14170 111796 14172
rect 111820 14170 111876 14172
rect 111900 14170 111956 14172
rect 111980 14170 112036 14172
rect 111740 14118 111786 14170
rect 111786 14118 111796 14170
rect 111820 14118 111850 14170
rect 111850 14118 111862 14170
rect 111862 14118 111876 14170
rect 111900 14118 111914 14170
rect 111914 14118 111926 14170
rect 111926 14118 111956 14170
rect 111980 14118 111990 14170
rect 111990 14118 112036 14170
rect 111740 14116 111796 14118
rect 111820 14116 111876 14118
rect 111900 14116 111956 14118
rect 111980 14116 112036 14118
rect 111740 13082 111796 13084
rect 111820 13082 111876 13084
rect 111900 13082 111956 13084
rect 111980 13082 112036 13084
rect 111740 13030 111786 13082
rect 111786 13030 111796 13082
rect 111820 13030 111850 13082
rect 111850 13030 111862 13082
rect 111862 13030 111876 13082
rect 111900 13030 111914 13082
rect 111914 13030 111926 13082
rect 111926 13030 111956 13082
rect 111980 13030 111990 13082
rect 111990 13030 112036 13082
rect 111740 13028 111796 13030
rect 111820 13028 111876 13030
rect 111900 13028 111956 13030
rect 111980 13028 112036 13030
rect 111740 11994 111796 11996
rect 111820 11994 111876 11996
rect 111900 11994 111956 11996
rect 111980 11994 112036 11996
rect 111740 11942 111786 11994
rect 111786 11942 111796 11994
rect 111820 11942 111850 11994
rect 111850 11942 111862 11994
rect 111862 11942 111876 11994
rect 111900 11942 111914 11994
rect 111914 11942 111926 11994
rect 111926 11942 111956 11994
rect 111980 11942 111990 11994
rect 111990 11942 112036 11994
rect 111740 11940 111796 11942
rect 111820 11940 111876 11942
rect 111900 11940 111956 11942
rect 111980 11940 112036 11942
rect 111740 10906 111796 10908
rect 111820 10906 111876 10908
rect 111900 10906 111956 10908
rect 111980 10906 112036 10908
rect 111740 10854 111786 10906
rect 111786 10854 111796 10906
rect 111820 10854 111850 10906
rect 111850 10854 111862 10906
rect 111862 10854 111876 10906
rect 111900 10854 111914 10906
rect 111914 10854 111926 10906
rect 111926 10854 111956 10906
rect 111980 10854 111990 10906
rect 111990 10854 112036 10906
rect 111740 10852 111796 10854
rect 111820 10852 111876 10854
rect 111900 10852 111956 10854
rect 111980 10852 112036 10854
rect 111740 9818 111796 9820
rect 111820 9818 111876 9820
rect 111900 9818 111956 9820
rect 111980 9818 112036 9820
rect 111740 9766 111786 9818
rect 111786 9766 111796 9818
rect 111820 9766 111850 9818
rect 111850 9766 111862 9818
rect 111862 9766 111876 9818
rect 111900 9766 111914 9818
rect 111914 9766 111926 9818
rect 111926 9766 111956 9818
rect 111980 9766 111990 9818
rect 111990 9766 112036 9818
rect 111740 9764 111796 9766
rect 111820 9764 111876 9766
rect 111900 9764 111956 9766
rect 111980 9764 112036 9766
rect 111740 8730 111796 8732
rect 111820 8730 111876 8732
rect 111900 8730 111956 8732
rect 111980 8730 112036 8732
rect 111740 8678 111786 8730
rect 111786 8678 111796 8730
rect 111820 8678 111850 8730
rect 111850 8678 111862 8730
rect 111862 8678 111876 8730
rect 111900 8678 111914 8730
rect 111914 8678 111926 8730
rect 111926 8678 111956 8730
rect 111980 8678 111990 8730
rect 111990 8678 112036 8730
rect 111740 8676 111796 8678
rect 111820 8676 111876 8678
rect 111900 8676 111956 8678
rect 111980 8676 112036 8678
rect 111740 7642 111796 7644
rect 111820 7642 111876 7644
rect 111900 7642 111956 7644
rect 111980 7642 112036 7644
rect 111740 7590 111786 7642
rect 111786 7590 111796 7642
rect 111820 7590 111850 7642
rect 111850 7590 111862 7642
rect 111862 7590 111876 7642
rect 111900 7590 111914 7642
rect 111914 7590 111926 7642
rect 111926 7590 111956 7642
rect 111980 7590 111990 7642
rect 111990 7590 112036 7642
rect 111740 7588 111796 7590
rect 111820 7588 111876 7590
rect 111900 7588 111956 7590
rect 111980 7588 112036 7590
rect 111740 6554 111796 6556
rect 111820 6554 111876 6556
rect 111900 6554 111956 6556
rect 111980 6554 112036 6556
rect 111740 6502 111786 6554
rect 111786 6502 111796 6554
rect 111820 6502 111850 6554
rect 111850 6502 111862 6554
rect 111862 6502 111876 6554
rect 111900 6502 111914 6554
rect 111914 6502 111926 6554
rect 111926 6502 111956 6554
rect 111980 6502 111990 6554
rect 111990 6502 112036 6554
rect 111740 6500 111796 6502
rect 111820 6500 111876 6502
rect 111900 6500 111956 6502
rect 111980 6500 112036 6502
rect 111740 5466 111796 5468
rect 111820 5466 111876 5468
rect 111900 5466 111956 5468
rect 111980 5466 112036 5468
rect 111740 5414 111786 5466
rect 111786 5414 111796 5466
rect 111820 5414 111850 5466
rect 111850 5414 111862 5466
rect 111862 5414 111876 5466
rect 111900 5414 111914 5466
rect 111914 5414 111926 5466
rect 111926 5414 111956 5466
rect 111980 5414 111990 5466
rect 111990 5414 112036 5466
rect 111740 5412 111796 5414
rect 111820 5412 111876 5414
rect 111900 5412 111956 5414
rect 111980 5412 112036 5414
rect 107290 3052 107346 3088
rect 107290 3032 107292 3052
rect 107292 3032 107344 3052
rect 107344 3032 107346 3052
rect 117226 12164 117282 12200
rect 117226 12144 117228 12164
rect 117228 12144 117280 12164
rect 117280 12144 117282 12164
rect 111740 4378 111796 4380
rect 111820 4378 111876 4380
rect 111900 4378 111956 4380
rect 111980 4378 112036 4380
rect 111740 4326 111786 4378
rect 111786 4326 111796 4378
rect 111820 4326 111850 4378
rect 111850 4326 111862 4378
rect 111862 4326 111876 4378
rect 111900 4326 111914 4378
rect 111914 4326 111926 4378
rect 111926 4326 111956 4378
rect 111980 4326 111990 4378
rect 111990 4326 112036 4378
rect 111740 4324 111796 4326
rect 111820 4324 111876 4326
rect 111900 4324 111956 4326
rect 111980 4324 112036 4326
rect 118054 34992 118110 35048
rect 118054 33496 118110 33552
rect 117962 29280 118018 29336
rect 118054 26424 118110 26480
rect 118054 23588 118110 23624
rect 118054 23568 118056 23588
rect 118056 23568 118108 23588
rect 118108 23568 118110 23588
rect 118054 22072 118110 22128
rect 117778 20712 117834 20768
rect 118054 19216 118110 19272
rect 117778 17856 117834 17912
rect 117778 15000 117834 15056
rect 117962 6432 118018 6488
rect 118054 4972 118056 4992
rect 118056 4972 118108 4992
rect 118108 4972 118110 4992
rect 118054 4936 118110 4972
rect 117962 3576 118018 3632
rect 111740 3290 111796 3292
rect 111820 3290 111876 3292
rect 111900 3290 111956 3292
rect 111980 3290 112036 3292
rect 111740 3238 111786 3290
rect 111786 3238 111796 3290
rect 111820 3238 111850 3290
rect 111850 3238 111862 3290
rect 111862 3238 111876 3290
rect 111900 3238 111914 3290
rect 111914 3238 111926 3290
rect 111926 3238 111956 3290
rect 111980 3238 111990 3290
rect 111990 3238 112036 3290
rect 111740 3236 111796 3238
rect 111820 3236 111876 3238
rect 111900 3236 111956 3238
rect 111980 3236 112036 3238
rect 110970 3032 111026 3088
rect 111740 2202 111796 2204
rect 111820 2202 111876 2204
rect 111900 2202 111956 2204
rect 111980 2202 112036 2204
rect 111740 2150 111786 2202
rect 111786 2150 111796 2202
rect 111820 2150 111850 2202
rect 111850 2150 111862 2202
rect 111862 2150 111876 2202
rect 111900 2150 111914 2202
rect 111914 2150 111926 2202
rect 111926 2150 111956 2202
rect 111980 2150 111990 2202
rect 111990 2150 112036 2202
rect 111740 2148 111796 2150
rect 111820 2148 111876 2150
rect 111900 2148 111956 2150
rect 111980 2148 112036 2150
rect 117962 2080 118018 2136
rect 118146 720 118202 776
<< metal3 >>
rect 117221 39266 117287 39269
rect 119200 39266 120000 39296
rect 117221 39264 120000 39266
rect 117221 39208 117226 39264
rect 117282 39208 120000 39264
rect 117221 39206 120000 39208
rect 117221 39203 117287 39206
rect 119200 39176 120000 39206
rect 0 39130 800 39160
rect 2773 39130 2839 39133
rect 0 39128 2839 39130
rect 0 39072 2778 39128
rect 2834 39072 2839 39128
rect 0 39070 2839 39072
rect 0 39040 800 39070
rect 2773 39067 2839 39070
rect 119200 37816 120000 37936
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 96370 37568 96686 37569
rect 96370 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96686 37568
rect 96370 37503 96686 37504
rect 1577 37498 1643 37501
rect 0 37496 1643 37498
rect 0 37440 1582 37496
rect 1638 37440 1643 37496
rect 0 37438 1643 37440
rect 0 37408 800 37438
rect 1577 37435 1643 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 81010 37024 81326 37025
rect 81010 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81326 37024
rect 81010 36959 81326 36960
rect 111730 37024 112046 37025
rect 111730 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112046 37024
rect 111730 36959 112046 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 96370 36480 96686 36481
rect 96370 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96686 36480
rect 96370 36415 96686 36416
rect 119200 36320 120000 36440
rect 19570 35936 19886 35937
rect 0 35866 800 35896
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 81010 35936 81326 35937
rect 81010 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81326 35936
rect 81010 35871 81326 35872
rect 111730 35936 112046 35937
rect 111730 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112046 35936
rect 111730 35871 112046 35872
rect 1485 35866 1551 35869
rect 0 35864 1551 35866
rect 0 35808 1490 35864
rect 1546 35808 1551 35864
rect 0 35806 1551 35808
rect 0 35776 800 35806
rect 1485 35803 1551 35806
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 96370 35392 96686 35393
rect 96370 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96686 35392
rect 96370 35327 96686 35328
rect 118049 35050 118115 35053
rect 119200 35050 120000 35080
rect 118049 35048 120000 35050
rect 118049 34992 118054 35048
rect 118110 34992 120000 35048
rect 118049 34990 120000 34992
rect 118049 34987 118115 34990
rect 119200 34960 120000 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 81010 34848 81326 34849
rect 81010 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81326 34848
rect 81010 34783 81326 34784
rect 111730 34848 112046 34849
rect 111730 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112046 34848
rect 111730 34783 112046 34784
rect 4210 34304 4526 34305
rect 0 34234 800 34264
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 96370 34304 96686 34305
rect 96370 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96686 34304
rect 96370 34239 96686 34240
rect 1577 34234 1643 34237
rect 0 34232 1643 34234
rect 0 34176 1582 34232
rect 1638 34176 1643 34232
rect 0 34174 1643 34176
rect 0 34144 800 34174
rect 1577 34171 1643 34174
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 81010 33760 81326 33761
rect 81010 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81326 33760
rect 81010 33695 81326 33696
rect 111730 33760 112046 33761
rect 111730 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112046 33760
rect 111730 33695 112046 33696
rect 118049 33554 118115 33557
rect 119200 33554 120000 33584
rect 118049 33552 120000 33554
rect 118049 33496 118054 33552
rect 118110 33496 120000 33552
rect 118049 33494 120000 33496
rect 118049 33491 118115 33494
rect 119200 33464 120000 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 96370 33216 96686 33217
rect 96370 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96686 33216
rect 96370 33151 96686 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 81010 32672 81326 32673
rect 81010 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81326 32672
rect 81010 32607 81326 32608
rect 111730 32672 112046 32673
rect 111730 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112046 32672
rect 111730 32607 112046 32608
rect 0 32466 800 32496
rect 1577 32466 1643 32469
rect 0 32464 1643 32466
rect 0 32408 1582 32464
rect 1638 32408 1643 32464
rect 0 32406 1643 32408
rect 0 32376 800 32406
rect 1577 32403 1643 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 96370 32128 96686 32129
rect 96370 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96686 32128
rect 119200 32104 120000 32224
rect 96370 32063 96686 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 81010 31584 81326 31585
rect 81010 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81326 31584
rect 81010 31519 81326 31520
rect 111730 31584 112046 31585
rect 111730 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112046 31584
rect 111730 31519 112046 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 96370 31040 96686 31041
rect 96370 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96686 31040
rect 96370 30975 96686 30976
rect 0 30744 800 30864
rect 119200 30608 120000 30728
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 81010 30496 81326 30497
rect 81010 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81326 30496
rect 81010 30431 81326 30432
rect 111730 30496 112046 30497
rect 111730 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112046 30496
rect 111730 30431 112046 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 96370 29952 96686 29953
rect 96370 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96686 29952
rect 96370 29887 96686 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 81010 29408 81326 29409
rect 81010 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81326 29408
rect 81010 29343 81326 29344
rect 111730 29408 112046 29409
rect 111730 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112046 29408
rect 111730 29343 112046 29344
rect 117957 29338 118023 29341
rect 119200 29338 120000 29368
rect 117957 29336 120000 29338
rect 117957 29280 117962 29336
rect 118018 29280 120000 29336
rect 117957 29278 120000 29280
rect 117957 29275 118023 29278
rect 119200 29248 120000 29278
rect 0 29202 800 29232
rect 1577 29202 1643 29205
rect 0 29200 1643 29202
rect 0 29144 1582 29200
rect 1638 29144 1643 29200
rect 0 29142 1643 29144
rect 0 29112 800 29142
rect 1577 29139 1643 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 96370 28864 96686 28865
rect 96370 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96686 28864
rect 96370 28799 96686 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 81010 28320 81326 28321
rect 81010 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81326 28320
rect 81010 28255 81326 28256
rect 111730 28320 112046 28321
rect 111730 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112046 28320
rect 111730 28255 112046 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 96370 27776 96686 27777
rect 96370 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96686 27776
rect 119200 27752 120000 27872
rect 96370 27711 96686 27712
rect 0 27480 800 27600
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 81010 27232 81326 27233
rect 81010 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81326 27232
rect 81010 27167 81326 27168
rect 111730 27232 112046 27233
rect 111730 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112046 27232
rect 111730 27167 112046 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 96370 26688 96686 26689
rect 96370 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96686 26688
rect 96370 26623 96686 26624
rect 118049 26482 118115 26485
rect 119200 26482 120000 26512
rect 118049 26480 120000 26482
rect 118049 26424 118054 26480
rect 118110 26424 120000 26480
rect 118049 26422 120000 26424
rect 118049 26419 118115 26422
rect 119200 26392 120000 26422
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 81010 26144 81326 26145
rect 81010 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81326 26144
rect 81010 26079 81326 26080
rect 111730 26144 112046 26145
rect 111730 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112046 26144
rect 111730 26079 112046 26080
rect 0 25802 800 25832
rect 1393 25802 1459 25805
rect 0 25800 1459 25802
rect 0 25744 1398 25800
rect 1454 25744 1459 25800
rect 0 25742 1459 25744
rect 0 25712 800 25742
rect 1393 25739 1459 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 96370 25600 96686 25601
rect 96370 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96686 25600
rect 96370 25535 96686 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 81010 25056 81326 25057
rect 81010 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81326 25056
rect 81010 24991 81326 24992
rect 111730 25056 112046 25057
rect 111730 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112046 25056
rect 111730 24991 112046 24992
rect 119200 24896 120000 25016
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 96370 24512 96686 24513
rect 96370 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96686 24512
rect 96370 24447 96686 24448
rect 0 24170 800 24200
rect 1577 24170 1643 24173
rect 0 24168 1643 24170
rect 0 24112 1582 24168
rect 1638 24112 1643 24168
rect 0 24110 1643 24112
rect 0 24080 800 24110
rect 1577 24107 1643 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 81010 23968 81326 23969
rect 81010 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81326 23968
rect 81010 23903 81326 23904
rect 111730 23968 112046 23969
rect 111730 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112046 23968
rect 111730 23903 112046 23904
rect 118049 23626 118115 23629
rect 119200 23626 120000 23656
rect 118049 23624 120000 23626
rect 118049 23568 118054 23624
rect 118110 23568 120000 23624
rect 118049 23566 120000 23568
rect 118049 23563 118115 23566
rect 119200 23536 120000 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 96370 23424 96686 23425
rect 96370 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96686 23424
rect 96370 23359 96686 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 81010 22880 81326 22881
rect 81010 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81326 22880
rect 81010 22815 81326 22816
rect 111730 22880 112046 22881
rect 111730 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112046 22880
rect 111730 22815 112046 22816
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 96370 22336 96686 22337
rect 96370 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96686 22336
rect 96370 22271 96686 22272
rect 118049 22130 118115 22133
rect 119200 22130 120000 22160
rect 118049 22128 120000 22130
rect 118049 22072 118054 22128
rect 118110 22072 120000 22128
rect 118049 22070 120000 22072
rect 118049 22067 118115 22070
rect 119200 22040 120000 22070
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 81010 21792 81326 21793
rect 81010 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81326 21792
rect 81010 21727 81326 21728
rect 111730 21792 112046 21793
rect 111730 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112046 21792
rect 111730 21727 112046 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 96370 21248 96686 21249
rect 96370 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96686 21248
rect 96370 21183 96686 21184
rect 0 20816 800 20936
rect 117773 20770 117839 20773
rect 119200 20770 120000 20800
rect 117773 20768 120000 20770
rect 117773 20712 117778 20768
rect 117834 20712 120000 20768
rect 117773 20710 120000 20712
rect 117773 20707 117839 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 81010 20704 81326 20705
rect 81010 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81326 20704
rect 81010 20639 81326 20640
rect 111730 20704 112046 20705
rect 111730 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112046 20704
rect 119200 20680 120000 20710
rect 111730 20639 112046 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 96370 20160 96686 20161
rect 96370 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96686 20160
rect 96370 20095 96686 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 81010 19616 81326 19617
rect 81010 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81326 19616
rect 81010 19551 81326 19552
rect 111730 19616 112046 19617
rect 111730 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112046 19616
rect 111730 19551 112046 19552
rect 118049 19274 118115 19277
rect 119200 19274 120000 19304
rect 118049 19272 120000 19274
rect 118049 19216 118054 19272
rect 118110 19216 120000 19272
rect 118049 19214 120000 19216
rect 118049 19211 118115 19214
rect 119200 19184 120000 19214
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 96370 19072 96686 19073
rect 96370 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96686 19072
rect 96370 19007 96686 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 81010 18528 81326 18529
rect 81010 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81326 18528
rect 81010 18463 81326 18464
rect 111730 18528 112046 18529
rect 111730 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112046 18528
rect 111730 18463 112046 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 96370 17984 96686 17985
rect 96370 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96686 17984
rect 96370 17919 96686 17920
rect 117773 17914 117839 17917
rect 119200 17914 120000 17944
rect 117773 17912 120000 17914
rect 117773 17856 117778 17912
rect 117834 17856 120000 17912
rect 117773 17854 120000 17856
rect 117773 17851 117839 17854
rect 119200 17824 120000 17854
rect 0 17506 800 17536
rect 1393 17506 1459 17509
rect 0 17504 1459 17506
rect 0 17448 1398 17504
rect 1454 17448 1459 17504
rect 0 17446 1459 17448
rect 0 17416 800 17446
rect 1393 17443 1459 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 81010 17440 81326 17441
rect 81010 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81326 17440
rect 81010 17375 81326 17376
rect 111730 17440 112046 17441
rect 111730 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112046 17440
rect 111730 17375 112046 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 96370 16896 96686 16897
rect 96370 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96686 16896
rect 96370 16831 96686 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 81010 16352 81326 16353
rect 81010 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81326 16352
rect 81010 16287 81326 16288
rect 111730 16352 112046 16353
rect 111730 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112046 16352
rect 119200 16328 120000 16448
rect 111730 16287 112046 16288
rect 0 15784 800 15904
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 96370 15808 96686 15809
rect 96370 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96686 15808
rect 96370 15743 96686 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 81010 15264 81326 15265
rect 81010 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81326 15264
rect 81010 15199 81326 15200
rect 111730 15264 112046 15265
rect 111730 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112046 15264
rect 111730 15199 112046 15200
rect 117773 15058 117839 15061
rect 119200 15058 120000 15088
rect 117773 15056 120000 15058
rect 117773 15000 117778 15056
rect 117834 15000 120000 15056
rect 117773 14998 120000 15000
rect 117773 14995 117839 14998
rect 119200 14968 120000 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 96370 14720 96686 14721
rect 96370 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96686 14720
rect 96370 14655 96686 14656
rect 0 14242 800 14272
rect 1853 14242 1919 14245
rect 0 14240 1919 14242
rect 0 14184 1858 14240
rect 1914 14184 1919 14240
rect 0 14182 1919 14184
rect 0 14152 800 14182
rect 1853 14179 1919 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 81010 14176 81326 14177
rect 81010 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81326 14176
rect 81010 14111 81326 14112
rect 111730 14176 112046 14177
rect 111730 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112046 14176
rect 111730 14111 112046 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 96370 13632 96686 13633
rect 96370 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96686 13632
rect 96370 13567 96686 13568
rect 119200 13472 120000 13592
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 81010 13088 81326 13089
rect 81010 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81326 13088
rect 81010 13023 81326 13024
rect 111730 13088 112046 13089
rect 111730 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112046 13088
rect 111730 13023 112046 13024
rect 4210 12544 4526 12545
rect 0 12384 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 96370 12544 96686 12545
rect 96370 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96686 12544
rect 96370 12479 96686 12480
rect 117221 12202 117287 12205
rect 119200 12202 120000 12232
rect 117221 12200 120000 12202
rect 117221 12144 117226 12200
rect 117282 12144 120000 12200
rect 117221 12142 120000 12144
rect 117221 12139 117287 12142
rect 119200 12112 120000 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 81010 12000 81326 12001
rect 81010 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81326 12000
rect 81010 11935 81326 11936
rect 111730 12000 112046 12001
rect 111730 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112046 12000
rect 111730 11935 112046 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 96370 11456 96686 11457
rect 96370 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96686 11456
rect 96370 11391 96686 11392
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 81010 10912 81326 10913
rect 81010 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81326 10912
rect 81010 10847 81326 10848
rect 111730 10912 112046 10913
rect 111730 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112046 10912
rect 111730 10847 112046 10848
rect 1853 10842 1919 10845
rect 0 10840 1919 10842
rect 0 10784 1858 10840
rect 1914 10784 1919 10840
rect 0 10782 1919 10784
rect 0 10752 800 10782
rect 1853 10779 1919 10782
rect 119200 10616 120000 10736
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 96370 10368 96686 10369
rect 96370 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96686 10368
rect 96370 10303 96686 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 81010 9824 81326 9825
rect 81010 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81326 9824
rect 81010 9759 81326 9760
rect 111730 9824 112046 9825
rect 111730 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112046 9824
rect 111730 9759 112046 9760
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 96370 9280 96686 9281
rect 96370 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96686 9280
rect 119200 9256 120000 9376
rect 96370 9215 96686 9216
rect 1577 9210 1643 9213
rect 0 9208 1643 9210
rect 0 9152 1582 9208
rect 1638 9152 1643 9208
rect 0 9150 1643 9152
rect 0 9120 800 9150
rect 1577 9147 1643 9150
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 81010 8736 81326 8737
rect 81010 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81326 8736
rect 81010 8671 81326 8672
rect 111730 8736 112046 8737
rect 111730 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112046 8736
rect 111730 8671 112046 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 96370 8192 96686 8193
rect 96370 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96686 8192
rect 96370 8127 96686 8128
rect 119200 7760 120000 7880
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 81010 7648 81326 7649
rect 81010 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81326 7648
rect 81010 7583 81326 7584
rect 111730 7648 112046 7649
rect 111730 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112046 7648
rect 111730 7583 112046 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 96370 7104 96686 7105
rect 96370 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96686 7104
rect 96370 7039 96686 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 81010 6560 81326 6561
rect 81010 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81326 6560
rect 81010 6495 81326 6496
rect 111730 6560 112046 6561
rect 111730 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112046 6560
rect 111730 6495 112046 6496
rect 117957 6490 118023 6493
rect 119200 6490 120000 6520
rect 117957 6488 120000 6490
rect 117957 6432 117962 6488
rect 118018 6432 120000 6488
rect 117957 6430 120000 6432
rect 117957 6427 118023 6430
rect 119200 6400 120000 6430
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 96370 6016 96686 6017
rect 96370 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96686 6016
rect 96370 5951 96686 5952
rect 0 5720 800 5840
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 81010 5472 81326 5473
rect 81010 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81326 5472
rect 81010 5407 81326 5408
rect 111730 5472 112046 5473
rect 111730 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112046 5472
rect 111730 5407 112046 5408
rect 118049 4994 118115 4997
rect 119200 4994 120000 5024
rect 118049 4992 120000 4994
rect 118049 4936 118054 4992
rect 118110 4936 120000 4992
rect 118049 4934 120000 4936
rect 118049 4931 118115 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 96370 4928 96686 4929
rect 96370 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96686 4928
rect 119200 4904 120000 4934
rect 96370 4863 96686 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 81010 4384 81326 4385
rect 81010 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81326 4384
rect 81010 4319 81326 4320
rect 111730 4384 112046 4385
rect 111730 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112046 4384
rect 111730 4319 112046 4320
rect 0 4088 800 4208
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 96370 3840 96686 3841
rect 96370 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96686 3840
rect 96370 3775 96686 3776
rect 117957 3634 118023 3637
rect 119200 3634 120000 3664
rect 117957 3632 120000 3634
rect 117957 3576 117962 3632
rect 118018 3576 120000 3632
rect 117957 3574 120000 3576
rect 117957 3571 118023 3574
rect 119200 3544 120000 3574
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 81010 3296 81326 3297
rect 81010 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81326 3296
rect 81010 3231 81326 3232
rect 111730 3296 112046 3297
rect 111730 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112046 3296
rect 111730 3231 112046 3232
rect 107285 3090 107351 3093
rect 110965 3090 111031 3093
rect 107285 3088 111031 3090
rect 107285 3032 107290 3088
rect 107346 3032 110970 3088
rect 111026 3032 111031 3088
rect 107285 3030 111031 3032
rect 107285 3027 107351 3030
rect 110965 3027 111031 3030
rect 39665 2954 39731 2957
rect 47577 2954 47643 2957
rect 39665 2952 47643 2954
rect 39665 2896 39670 2952
rect 39726 2896 47582 2952
rect 47638 2896 47643 2952
rect 39665 2894 47643 2896
rect 39665 2891 39731 2894
rect 47577 2891 47643 2894
rect 50613 2954 50679 2957
rect 104249 2954 104315 2957
rect 50613 2952 104315 2954
rect 50613 2896 50618 2952
rect 50674 2896 104254 2952
rect 104310 2896 104315 2952
rect 50613 2894 104315 2896
rect 50613 2891 50679 2894
rect 104249 2891 104315 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 96370 2752 96686 2753
rect 96370 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96686 2752
rect 96370 2687 96686 2688
rect 0 2456 800 2576
rect 62665 2410 62731 2413
rect 65701 2410 65767 2413
rect 62665 2408 65767 2410
rect 62665 2352 62670 2408
rect 62726 2352 65706 2408
rect 65762 2352 65767 2408
rect 62665 2350 65767 2352
rect 62665 2347 62731 2350
rect 65701 2347 65767 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 81010 2208 81326 2209
rect 81010 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81326 2208
rect 81010 2143 81326 2144
rect 111730 2208 112046 2209
rect 111730 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112046 2208
rect 111730 2143 112046 2144
rect 117957 2138 118023 2141
rect 119200 2138 120000 2168
rect 117957 2136 120000 2138
rect 117957 2080 117962 2136
rect 118018 2080 120000 2136
rect 117957 2078 120000 2080
rect 117957 2075 118023 2078
rect 119200 2048 120000 2078
rect 0 914 800 944
rect 1393 914 1459 917
rect 0 912 1459 914
rect 0 856 1398 912
rect 1454 856 1459 912
rect 0 854 1459 856
rect 0 824 800 854
rect 1393 851 1459 854
rect 118141 778 118207 781
rect 119200 778 120000 808
rect 118141 776 120000 778
rect 118141 720 118146 776
rect 118202 720 120000 776
rect 118141 718 120000 720
rect 118141 715 118207 718
rect 119200 688 120000 718
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 96376 37564 96440 37568
rect 96376 37508 96380 37564
rect 96380 37508 96436 37564
rect 96436 37508 96440 37564
rect 96376 37504 96440 37508
rect 96456 37564 96520 37568
rect 96456 37508 96460 37564
rect 96460 37508 96516 37564
rect 96516 37508 96520 37564
rect 96456 37504 96520 37508
rect 96536 37564 96600 37568
rect 96536 37508 96540 37564
rect 96540 37508 96596 37564
rect 96596 37508 96600 37564
rect 96536 37504 96600 37508
rect 96616 37564 96680 37568
rect 96616 37508 96620 37564
rect 96620 37508 96676 37564
rect 96676 37508 96680 37564
rect 96616 37504 96680 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 81016 37020 81080 37024
rect 81016 36964 81020 37020
rect 81020 36964 81076 37020
rect 81076 36964 81080 37020
rect 81016 36960 81080 36964
rect 81096 37020 81160 37024
rect 81096 36964 81100 37020
rect 81100 36964 81156 37020
rect 81156 36964 81160 37020
rect 81096 36960 81160 36964
rect 81176 37020 81240 37024
rect 81176 36964 81180 37020
rect 81180 36964 81236 37020
rect 81236 36964 81240 37020
rect 81176 36960 81240 36964
rect 81256 37020 81320 37024
rect 81256 36964 81260 37020
rect 81260 36964 81316 37020
rect 81316 36964 81320 37020
rect 81256 36960 81320 36964
rect 111736 37020 111800 37024
rect 111736 36964 111740 37020
rect 111740 36964 111796 37020
rect 111796 36964 111800 37020
rect 111736 36960 111800 36964
rect 111816 37020 111880 37024
rect 111816 36964 111820 37020
rect 111820 36964 111876 37020
rect 111876 36964 111880 37020
rect 111816 36960 111880 36964
rect 111896 37020 111960 37024
rect 111896 36964 111900 37020
rect 111900 36964 111956 37020
rect 111956 36964 111960 37020
rect 111896 36960 111960 36964
rect 111976 37020 112040 37024
rect 111976 36964 111980 37020
rect 111980 36964 112036 37020
rect 112036 36964 112040 37020
rect 111976 36960 112040 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 96376 36476 96440 36480
rect 96376 36420 96380 36476
rect 96380 36420 96436 36476
rect 96436 36420 96440 36476
rect 96376 36416 96440 36420
rect 96456 36476 96520 36480
rect 96456 36420 96460 36476
rect 96460 36420 96516 36476
rect 96516 36420 96520 36476
rect 96456 36416 96520 36420
rect 96536 36476 96600 36480
rect 96536 36420 96540 36476
rect 96540 36420 96596 36476
rect 96596 36420 96600 36476
rect 96536 36416 96600 36420
rect 96616 36476 96680 36480
rect 96616 36420 96620 36476
rect 96620 36420 96676 36476
rect 96676 36420 96680 36476
rect 96616 36416 96680 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 81016 35932 81080 35936
rect 81016 35876 81020 35932
rect 81020 35876 81076 35932
rect 81076 35876 81080 35932
rect 81016 35872 81080 35876
rect 81096 35932 81160 35936
rect 81096 35876 81100 35932
rect 81100 35876 81156 35932
rect 81156 35876 81160 35932
rect 81096 35872 81160 35876
rect 81176 35932 81240 35936
rect 81176 35876 81180 35932
rect 81180 35876 81236 35932
rect 81236 35876 81240 35932
rect 81176 35872 81240 35876
rect 81256 35932 81320 35936
rect 81256 35876 81260 35932
rect 81260 35876 81316 35932
rect 81316 35876 81320 35932
rect 81256 35872 81320 35876
rect 111736 35932 111800 35936
rect 111736 35876 111740 35932
rect 111740 35876 111796 35932
rect 111796 35876 111800 35932
rect 111736 35872 111800 35876
rect 111816 35932 111880 35936
rect 111816 35876 111820 35932
rect 111820 35876 111876 35932
rect 111876 35876 111880 35932
rect 111816 35872 111880 35876
rect 111896 35932 111960 35936
rect 111896 35876 111900 35932
rect 111900 35876 111956 35932
rect 111956 35876 111960 35932
rect 111896 35872 111960 35876
rect 111976 35932 112040 35936
rect 111976 35876 111980 35932
rect 111980 35876 112036 35932
rect 112036 35876 112040 35932
rect 111976 35872 112040 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 96376 35388 96440 35392
rect 96376 35332 96380 35388
rect 96380 35332 96436 35388
rect 96436 35332 96440 35388
rect 96376 35328 96440 35332
rect 96456 35388 96520 35392
rect 96456 35332 96460 35388
rect 96460 35332 96516 35388
rect 96516 35332 96520 35388
rect 96456 35328 96520 35332
rect 96536 35388 96600 35392
rect 96536 35332 96540 35388
rect 96540 35332 96596 35388
rect 96596 35332 96600 35388
rect 96536 35328 96600 35332
rect 96616 35388 96680 35392
rect 96616 35332 96620 35388
rect 96620 35332 96676 35388
rect 96676 35332 96680 35388
rect 96616 35328 96680 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 81016 34844 81080 34848
rect 81016 34788 81020 34844
rect 81020 34788 81076 34844
rect 81076 34788 81080 34844
rect 81016 34784 81080 34788
rect 81096 34844 81160 34848
rect 81096 34788 81100 34844
rect 81100 34788 81156 34844
rect 81156 34788 81160 34844
rect 81096 34784 81160 34788
rect 81176 34844 81240 34848
rect 81176 34788 81180 34844
rect 81180 34788 81236 34844
rect 81236 34788 81240 34844
rect 81176 34784 81240 34788
rect 81256 34844 81320 34848
rect 81256 34788 81260 34844
rect 81260 34788 81316 34844
rect 81316 34788 81320 34844
rect 81256 34784 81320 34788
rect 111736 34844 111800 34848
rect 111736 34788 111740 34844
rect 111740 34788 111796 34844
rect 111796 34788 111800 34844
rect 111736 34784 111800 34788
rect 111816 34844 111880 34848
rect 111816 34788 111820 34844
rect 111820 34788 111876 34844
rect 111876 34788 111880 34844
rect 111816 34784 111880 34788
rect 111896 34844 111960 34848
rect 111896 34788 111900 34844
rect 111900 34788 111956 34844
rect 111956 34788 111960 34844
rect 111896 34784 111960 34788
rect 111976 34844 112040 34848
rect 111976 34788 111980 34844
rect 111980 34788 112036 34844
rect 112036 34788 112040 34844
rect 111976 34784 112040 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 96376 34300 96440 34304
rect 96376 34244 96380 34300
rect 96380 34244 96436 34300
rect 96436 34244 96440 34300
rect 96376 34240 96440 34244
rect 96456 34300 96520 34304
rect 96456 34244 96460 34300
rect 96460 34244 96516 34300
rect 96516 34244 96520 34300
rect 96456 34240 96520 34244
rect 96536 34300 96600 34304
rect 96536 34244 96540 34300
rect 96540 34244 96596 34300
rect 96596 34244 96600 34300
rect 96536 34240 96600 34244
rect 96616 34300 96680 34304
rect 96616 34244 96620 34300
rect 96620 34244 96676 34300
rect 96676 34244 96680 34300
rect 96616 34240 96680 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 81016 33756 81080 33760
rect 81016 33700 81020 33756
rect 81020 33700 81076 33756
rect 81076 33700 81080 33756
rect 81016 33696 81080 33700
rect 81096 33756 81160 33760
rect 81096 33700 81100 33756
rect 81100 33700 81156 33756
rect 81156 33700 81160 33756
rect 81096 33696 81160 33700
rect 81176 33756 81240 33760
rect 81176 33700 81180 33756
rect 81180 33700 81236 33756
rect 81236 33700 81240 33756
rect 81176 33696 81240 33700
rect 81256 33756 81320 33760
rect 81256 33700 81260 33756
rect 81260 33700 81316 33756
rect 81316 33700 81320 33756
rect 81256 33696 81320 33700
rect 111736 33756 111800 33760
rect 111736 33700 111740 33756
rect 111740 33700 111796 33756
rect 111796 33700 111800 33756
rect 111736 33696 111800 33700
rect 111816 33756 111880 33760
rect 111816 33700 111820 33756
rect 111820 33700 111876 33756
rect 111876 33700 111880 33756
rect 111816 33696 111880 33700
rect 111896 33756 111960 33760
rect 111896 33700 111900 33756
rect 111900 33700 111956 33756
rect 111956 33700 111960 33756
rect 111896 33696 111960 33700
rect 111976 33756 112040 33760
rect 111976 33700 111980 33756
rect 111980 33700 112036 33756
rect 112036 33700 112040 33756
rect 111976 33696 112040 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 96376 33212 96440 33216
rect 96376 33156 96380 33212
rect 96380 33156 96436 33212
rect 96436 33156 96440 33212
rect 96376 33152 96440 33156
rect 96456 33212 96520 33216
rect 96456 33156 96460 33212
rect 96460 33156 96516 33212
rect 96516 33156 96520 33212
rect 96456 33152 96520 33156
rect 96536 33212 96600 33216
rect 96536 33156 96540 33212
rect 96540 33156 96596 33212
rect 96596 33156 96600 33212
rect 96536 33152 96600 33156
rect 96616 33212 96680 33216
rect 96616 33156 96620 33212
rect 96620 33156 96676 33212
rect 96676 33156 96680 33212
rect 96616 33152 96680 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 81016 32668 81080 32672
rect 81016 32612 81020 32668
rect 81020 32612 81076 32668
rect 81076 32612 81080 32668
rect 81016 32608 81080 32612
rect 81096 32668 81160 32672
rect 81096 32612 81100 32668
rect 81100 32612 81156 32668
rect 81156 32612 81160 32668
rect 81096 32608 81160 32612
rect 81176 32668 81240 32672
rect 81176 32612 81180 32668
rect 81180 32612 81236 32668
rect 81236 32612 81240 32668
rect 81176 32608 81240 32612
rect 81256 32668 81320 32672
rect 81256 32612 81260 32668
rect 81260 32612 81316 32668
rect 81316 32612 81320 32668
rect 81256 32608 81320 32612
rect 111736 32668 111800 32672
rect 111736 32612 111740 32668
rect 111740 32612 111796 32668
rect 111796 32612 111800 32668
rect 111736 32608 111800 32612
rect 111816 32668 111880 32672
rect 111816 32612 111820 32668
rect 111820 32612 111876 32668
rect 111876 32612 111880 32668
rect 111816 32608 111880 32612
rect 111896 32668 111960 32672
rect 111896 32612 111900 32668
rect 111900 32612 111956 32668
rect 111956 32612 111960 32668
rect 111896 32608 111960 32612
rect 111976 32668 112040 32672
rect 111976 32612 111980 32668
rect 111980 32612 112036 32668
rect 112036 32612 112040 32668
rect 111976 32608 112040 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 96376 32124 96440 32128
rect 96376 32068 96380 32124
rect 96380 32068 96436 32124
rect 96436 32068 96440 32124
rect 96376 32064 96440 32068
rect 96456 32124 96520 32128
rect 96456 32068 96460 32124
rect 96460 32068 96516 32124
rect 96516 32068 96520 32124
rect 96456 32064 96520 32068
rect 96536 32124 96600 32128
rect 96536 32068 96540 32124
rect 96540 32068 96596 32124
rect 96596 32068 96600 32124
rect 96536 32064 96600 32068
rect 96616 32124 96680 32128
rect 96616 32068 96620 32124
rect 96620 32068 96676 32124
rect 96676 32068 96680 32124
rect 96616 32064 96680 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 81016 31580 81080 31584
rect 81016 31524 81020 31580
rect 81020 31524 81076 31580
rect 81076 31524 81080 31580
rect 81016 31520 81080 31524
rect 81096 31580 81160 31584
rect 81096 31524 81100 31580
rect 81100 31524 81156 31580
rect 81156 31524 81160 31580
rect 81096 31520 81160 31524
rect 81176 31580 81240 31584
rect 81176 31524 81180 31580
rect 81180 31524 81236 31580
rect 81236 31524 81240 31580
rect 81176 31520 81240 31524
rect 81256 31580 81320 31584
rect 81256 31524 81260 31580
rect 81260 31524 81316 31580
rect 81316 31524 81320 31580
rect 81256 31520 81320 31524
rect 111736 31580 111800 31584
rect 111736 31524 111740 31580
rect 111740 31524 111796 31580
rect 111796 31524 111800 31580
rect 111736 31520 111800 31524
rect 111816 31580 111880 31584
rect 111816 31524 111820 31580
rect 111820 31524 111876 31580
rect 111876 31524 111880 31580
rect 111816 31520 111880 31524
rect 111896 31580 111960 31584
rect 111896 31524 111900 31580
rect 111900 31524 111956 31580
rect 111956 31524 111960 31580
rect 111896 31520 111960 31524
rect 111976 31580 112040 31584
rect 111976 31524 111980 31580
rect 111980 31524 112036 31580
rect 112036 31524 112040 31580
rect 111976 31520 112040 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 96376 31036 96440 31040
rect 96376 30980 96380 31036
rect 96380 30980 96436 31036
rect 96436 30980 96440 31036
rect 96376 30976 96440 30980
rect 96456 31036 96520 31040
rect 96456 30980 96460 31036
rect 96460 30980 96516 31036
rect 96516 30980 96520 31036
rect 96456 30976 96520 30980
rect 96536 31036 96600 31040
rect 96536 30980 96540 31036
rect 96540 30980 96596 31036
rect 96596 30980 96600 31036
rect 96536 30976 96600 30980
rect 96616 31036 96680 31040
rect 96616 30980 96620 31036
rect 96620 30980 96676 31036
rect 96676 30980 96680 31036
rect 96616 30976 96680 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 81016 30492 81080 30496
rect 81016 30436 81020 30492
rect 81020 30436 81076 30492
rect 81076 30436 81080 30492
rect 81016 30432 81080 30436
rect 81096 30492 81160 30496
rect 81096 30436 81100 30492
rect 81100 30436 81156 30492
rect 81156 30436 81160 30492
rect 81096 30432 81160 30436
rect 81176 30492 81240 30496
rect 81176 30436 81180 30492
rect 81180 30436 81236 30492
rect 81236 30436 81240 30492
rect 81176 30432 81240 30436
rect 81256 30492 81320 30496
rect 81256 30436 81260 30492
rect 81260 30436 81316 30492
rect 81316 30436 81320 30492
rect 81256 30432 81320 30436
rect 111736 30492 111800 30496
rect 111736 30436 111740 30492
rect 111740 30436 111796 30492
rect 111796 30436 111800 30492
rect 111736 30432 111800 30436
rect 111816 30492 111880 30496
rect 111816 30436 111820 30492
rect 111820 30436 111876 30492
rect 111876 30436 111880 30492
rect 111816 30432 111880 30436
rect 111896 30492 111960 30496
rect 111896 30436 111900 30492
rect 111900 30436 111956 30492
rect 111956 30436 111960 30492
rect 111896 30432 111960 30436
rect 111976 30492 112040 30496
rect 111976 30436 111980 30492
rect 111980 30436 112036 30492
rect 112036 30436 112040 30492
rect 111976 30432 112040 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 96376 29948 96440 29952
rect 96376 29892 96380 29948
rect 96380 29892 96436 29948
rect 96436 29892 96440 29948
rect 96376 29888 96440 29892
rect 96456 29948 96520 29952
rect 96456 29892 96460 29948
rect 96460 29892 96516 29948
rect 96516 29892 96520 29948
rect 96456 29888 96520 29892
rect 96536 29948 96600 29952
rect 96536 29892 96540 29948
rect 96540 29892 96596 29948
rect 96596 29892 96600 29948
rect 96536 29888 96600 29892
rect 96616 29948 96680 29952
rect 96616 29892 96620 29948
rect 96620 29892 96676 29948
rect 96676 29892 96680 29948
rect 96616 29888 96680 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 81016 29404 81080 29408
rect 81016 29348 81020 29404
rect 81020 29348 81076 29404
rect 81076 29348 81080 29404
rect 81016 29344 81080 29348
rect 81096 29404 81160 29408
rect 81096 29348 81100 29404
rect 81100 29348 81156 29404
rect 81156 29348 81160 29404
rect 81096 29344 81160 29348
rect 81176 29404 81240 29408
rect 81176 29348 81180 29404
rect 81180 29348 81236 29404
rect 81236 29348 81240 29404
rect 81176 29344 81240 29348
rect 81256 29404 81320 29408
rect 81256 29348 81260 29404
rect 81260 29348 81316 29404
rect 81316 29348 81320 29404
rect 81256 29344 81320 29348
rect 111736 29404 111800 29408
rect 111736 29348 111740 29404
rect 111740 29348 111796 29404
rect 111796 29348 111800 29404
rect 111736 29344 111800 29348
rect 111816 29404 111880 29408
rect 111816 29348 111820 29404
rect 111820 29348 111876 29404
rect 111876 29348 111880 29404
rect 111816 29344 111880 29348
rect 111896 29404 111960 29408
rect 111896 29348 111900 29404
rect 111900 29348 111956 29404
rect 111956 29348 111960 29404
rect 111896 29344 111960 29348
rect 111976 29404 112040 29408
rect 111976 29348 111980 29404
rect 111980 29348 112036 29404
rect 112036 29348 112040 29404
rect 111976 29344 112040 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 96376 28860 96440 28864
rect 96376 28804 96380 28860
rect 96380 28804 96436 28860
rect 96436 28804 96440 28860
rect 96376 28800 96440 28804
rect 96456 28860 96520 28864
rect 96456 28804 96460 28860
rect 96460 28804 96516 28860
rect 96516 28804 96520 28860
rect 96456 28800 96520 28804
rect 96536 28860 96600 28864
rect 96536 28804 96540 28860
rect 96540 28804 96596 28860
rect 96596 28804 96600 28860
rect 96536 28800 96600 28804
rect 96616 28860 96680 28864
rect 96616 28804 96620 28860
rect 96620 28804 96676 28860
rect 96676 28804 96680 28860
rect 96616 28800 96680 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 81016 28316 81080 28320
rect 81016 28260 81020 28316
rect 81020 28260 81076 28316
rect 81076 28260 81080 28316
rect 81016 28256 81080 28260
rect 81096 28316 81160 28320
rect 81096 28260 81100 28316
rect 81100 28260 81156 28316
rect 81156 28260 81160 28316
rect 81096 28256 81160 28260
rect 81176 28316 81240 28320
rect 81176 28260 81180 28316
rect 81180 28260 81236 28316
rect 81236 28260 81240 28316
rect 81176 28256 81240 28260
rect 81256 28316 81320 28320
rect 81256 28260 81260 28316
rect 81260 28260 81316 28316
rect 81316 28260 81320 28316
rect 81256 28256 81320 28260
rect 111736 28316 111800 28320
rect 111736 28260 111740 28316
rect 111740 28260 111796 28316
rect 111796 28260 111800 28316
rect 111736 28256 111800 28260
rect 111816 28316 111880 28320
rect 111816 28260 111820 28316
rect 111820 28260 111876 28316
rect 111876 28260 111880 28316
rect 111816 28256 111880 28260
rect 111896 28316 111960 28320
rect 111896 28260 111900 28316
rect 111900 28260 111956 28316
rect 111956 28260 111960 28316
rect 111896 28256 111960 28260
rect 111976 28316 112040 28320
rect 111976 28260 111980 28316
rect 111980 28260 112036 28316
rect 112036 28260 112040 28316
rect 111976 28256 112040 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 96376 27772 96440 27776
rect 96376 27716 96380 27772
rect 96380 27716 96436 27772
rect 96436 27716 96440 27772
rect 96376 27712 96440 27716
rect 96456 27772 96520 27776
rect 96456 27716 96460 27772
rect 96460 27716 96516 27772
rect 96516 27716 96520 27772
rect 96456 27712 96520 27716
rect 96536 27772 96600 27776
rect 96536 27716 96540 27772
rect 96540 27716 96596 27772
rect 96596 27716 96600 27772
rect 96536 27712 96600 27716
rect 96616 27772 96680 27776
rect 96616 27716 96620 27772
rect 96620 27716 96676 27772
rect 96676 27716 96680 27772
rect 96616 27712 96680 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 81016 27228 81080 27232
rect 81016 27172 81020 27228
rect 81020 27172 81076 27228
rect 81076 27172 81080 27228
rect 81016 27168 81080 27172
rect 81096 27228 81160 27232
rect 81096 27172 81100 27228
rect 81100 27172 81156 27228
rect 81156 27172 81160 27228
rect 81096 27168 81160 27172
rect 81176 27228 81240 27232
rect 81176 27172 81180 27228
rect 81180 27172 81236 27228
rect 81236 27172 81240 27228
rect 81176 27168 81240 27172
rect 81256 27228 81320 27232
rect 81256 27172 81260 27228
rect 81260 27172 81316 27228
rect 81316 27172 81320 27228
rect 81256 27168 81320 27172
rect 111736 27228 111800 27232
rect 111736 27172 111740 27228
rect 111740 27172 111796 27228
rect 111796 27172 111800 27228
rect 111736 27168 111800 27172
rect 111816 27228 111880 27232
rect 111816 27172 111820 27228
rect 111820 27172 111876 27228
rect 111876 27172 111880 27228
rect 111816 27168 111880 27172
rect 111896 27228 111960 27232
rect 111896 27172 111900 27228
rect 111900 27172 111956 27228
rect 111956 27172 111960 27228
rect 111896 27168 111960 27172
rect 111976 27228 112040 27232
rect 111976 27172 111980 27228
rect 111980 27172 112036 27228
rect 112036 27172 112040 27228
rect 111976 27168 112040 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 96376 26684 96440 26688
rect 96376 26628 96380 26684
rect 96380 26628 96436 26684
rect 96436 26628 96440 26684
rect 96376 26624 96440 26628
rect 96456 26684 96520 26688
rect 96456 26628 96460 26684
rect 96460 26628 96516 26684
rect 96516 26628 96520 26684
rect 96456 26624 96520 26628
rect 96536 26684 96600 26688
rect 96536 26628 96540 26684
rect 96540 26628 96596 26684
rect 96596 26628 96600 26684
rect 96536 26624 96600 26628
rect 96616 26684 96680 26688
rect 96616 26628 96620 26684
rect 96620 26628 96676 26684
rect 96676 26628 96680 26684
rect 96616 26624 96680 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 81016 26140 81080 26144
rect 81016 26084 81020 26140
rect 81020 26084 81076 26140
rect 81076 26084 81080 26140
rect 81016 26080 81080 26084
rect 81096 26140 81160 26144
rect 81096 26084 81100 26140
rect 81100 26084 81156 26140
rect 81156 26084 81160 26140
rect 81096 26080 81160 26084
rect 81176 26140 81240 26144
rect 81176 26084 81180 26140
rect 81180 26084 81236 26140
rect 81236 26084 81240 26140
rect 81176 26080 81240 26084
rect 81256 26140 81320 26144
rect 81256 26084 81260 26140
rect 81260 26084 81316 26140
rect 81316 26084 81320 26140
rect 81256 26080 81320 26084
rect 111736 26140 111800 26144
rect 111736 26084 111740 26140
rect 111740 26084 111796 26140
rect 111796 26084 111800 26140
rect 111736 26080 111800 26084
rect 111816 26140 111880 26144
rect 111816 26084 111820 26140
rect 111820 26084 111876 26140
rect 111876 26084 111880 26140
rect 111816 26080 111880 26084
rect 111896 26140 111960 26144
rect 111896 26084 111900 26140
rect 111900 26084 111956 26140
rect 111956 26084 111960 26140
rect 111896 26080 111960 26084
rect 111976 26140 112040 26144
rect 111976 26084 111980 26140
rect 111980 26084 112036 26140
rect 112036 26084 112040 26140
rect 111976 26080 112040 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 96376 25596 96440 25600
rect 96376 25540 96380 25596
rect 96380 25540 96436 25596
rect 96436 25540 96440 25596
rect 96376 25536 96440 25540
rect 96456 25596 96520 25600
rect 96456 25540 96460 25596
rect 96460 25540 96516 25596
rect 96516 25540 96520 25596
rect 96456 25536 96520 25540
rect 96536 25596 96600 25600
rect 96536 25540 96540 25596
rect 96540 25540 96596 25596
rect 96596 25540 96600 25596
rect 96536 25536 96600 25540
rect 96616 25596 96680 25600
rect 96616 25540 96620 25596
rect 96620 25540 96676 25596
rect 96676 25540 96680 25596
rect 96616 25536 96680 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 81016 25052 81080 25056
rect 81016 24996 81020 25052
rect 81020 24996 81076 25052
rect 81076 24996 81080 25052
rect 81016 24992 81080 24996
rect 81096 25052 81160 25056
rect 81096 24996 81100 25052
rect 81100 24996 81156 25052
rect 81156 24996 81160 25052
rect 81096 24992 81160 24996
rect 81176 25052 81240 25056
rect 81176 24996 81180 25052
rect 81180 24996 81236 25052
rect 81236 24996 81240 25052
rect 81176 24992 81240 24996
rect 81256 25052 81320 25056
rect 81256 24996 81260 25052
rect 81260 24996 81316 25052
rect 81316 24996 81320 25052
rect 81256 24992 81320 24996
rect 111736 25052 111800 25056
rect 111736 24996 111740 25052
rect 111740 24996 111796 25052
rect 111796 24996 111800 25052
rect 111736 24992 111800 24996
rect 111816 25052 111880 25056
rect 111816 24996 111820 25052
rect 111820 24996 111876 25052
rect 111876 24996 111880 25052
rect 111816 24992 111880 24996
rect 111896 25052 111960 25056
rect 111896 24996 111900 25052
rect 111900 24996 111956 25052
rect 111956 24996 111960 25052
rect 111896 24992 111960 24996
rect 111976 25052 112040 25056
rect 111976 24996 111980 25052
rect 111980 24996 112036 25052
rect 112036 24996 112040 25052
rect 111976 24992 112040 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 96376 24508 96440 24512
rect 96376 24452 96380 24508
rect 96380 24452 96436 24508
rect 96436 24452 96440 24508
rect 96376 24448 96440 24452
rect 96456 24508 96520 24512
rect 96456 24452 96460 24508
rect 96460 24452 96516 24508
rect 96516 24452 96520 24508
rect 96456 24448 96520 24452
rect 96536 24508 96600 24512
rect 96536 24452 96540 24508
rect 96540 24452 96596 24508
rect 96596 24452 96600 24508
rect 96536 24448 96600 24452
rect 96616 24508 96680 24512
rect 96616 24452 96620 24508
rect 96620 24452 96676 24508
rect 96676 24452 96680 24508
rect 96616 24448 96680 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 81016 23964 81080 23968
rect 81016 23908 81020 23964
rect 81020 23908 81076 23964
rect 81076 23908 81080 23964
rect 81016 23904 81080 23908
rect 81096 23964 81160 23968
rect 81096 23908 81100 23964
rect 81100 23908 81156 23964
rect 81156 23908 81160 23964
rect 81096 23904 81160 23908
rect 81176 23964 81240 23968
rect 81176 23908 81180 23964
rect 81180 23908 81236 23964
rect 81236 23908 81240 23964
rect 81176 23904 81240 23908
rect 81256 23964 81320 23968
rect 81256 23908 81260 23964
rect 81260 23908 81316 23964
rect 81316 23908 81320 23964
rect 81256 23904 81320 23908
rect 111736 23964 111800 23968
rect 111736 23908 111740 23964
rect 111740 23908 111796 23964
rect 111796 23908 111800 23964
rect 111736 23904 111800 23908
rect 111816 23964 111880 23968
rect 111816 23908 111820 23964
rect 111820 23908 111876 23964
rect 111876 23908 111880 23964
rect 111816 23904 111880 23908
rect 111896 23964 111960 23968
rect 111896 23908 111900 23964
rect 111900 23908 111956 23964
rect 111956 23908 111960 23964
rect 111896 23904 111960 23908
rect 111976 23964 112040 23968
rect 111976 23908 111980 23964
rect 111980 23908 112036 23964
rect 112036 23908 112040 23964
rect 111976 23904 112040 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 96376 23420 96440 23424
rect 96376 23364 96380 23420
rect 96380 23364 96436 23420
rect 96436 23364 96440 23420
rect 96376 23360 96440 23364
rect 96456 23420 96520 23424
rect 96456 23364 96460 23420
rect 96460 23364 96516 23420
rect 96516 23364 96520 23420
rect 96456 23360 96520 23364
rect 96536 23420 96600 23424
rect 96536 23364 96540 23420
rect 96540 23364 96596 23420
rect 96596 23364 96600 23420
rect 96536 23360 96600 23364
rect 96616 23420 96680 23424
rect 96616 23364 96620 23420
rect 96620 23364 96676 23420
rect 96676 23364 96680 23420
rect 96616 23360 96680 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 81016 22876 81080 22880
rect 81016 22820 81020 22876
rect 81020 22820 81076 22876
rect 81076 22820 81080 22876
rect 81016 22816 81080 22820
rect 81096 22876 81160 22880
rect 81096 22820 81100 22876
rect 81100 22820 81156 22876
rect 81156 22820 81160 22876
rect 81096 22816 81160 22820
rect 81176 22876 81240 22880
rect 81176 22820 81180 22876
rect 81180 22820 81236 22876
rect 81236 22820 81240 22876
rect 81176 22816 81240 22820
rect 81256 22876 81320 22880
rect 81256 22820 81260 22876
rect 81260 22820 81316 22876
rect 81316 22820 81320 22876
rect 81256 22816 81320 22820
rect 111736 22876 111800 22880
rect 111736 22820 111740 22876
rect 111740 22820 111796 22876
rect 111796 22820 111800 22876
rect 111736 22816 111800 22820
rect 111816 22876 111880 22880
rect 111816 22820 111820 22876
rect 111820 22820 111876 22876
rect 111876 22820 111880 22876
rect 111816 22816 111880 22820
rect 111896 22876 111960 22880
rect 111896 22820 111900 22876
rect 111900 22820 111956 22876
rect 111956 22820 111960 22876
rect 111896 22816 111960 22820
rect 111976 22876 112040 22880
rect 111976 22820 111980 22876
rect 111980 22820 112036 22876
rect 112036 22820 112040 22876
rect 111976 22816 112040 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 96376 22332 96440 22336
rect 96376 22276 96380 22332
rect 96380 22276 96436 22332
rect 96436 22276 96440 22332
rect 96376 22272 96440 22276
rect 96456 22332 96520 22336
rect 96456 22276 96460 22332
rect 96460 22276 96516 22332
rect 96516 22276 96520 22332
rect 96456 22272 96520 22276
rect 96536 22332 96600 22336
rect 96536 22276 96540 22332
rect 96540 22276 96596 22332
rect 96596 22276 96600 22332
rect 96536 22272 96600 22276
rect 96616 22332 96680 22336
rect 96616 22276 96620 22332
rect 96620 22276 96676 22332
rect 96676 22276 96680 22332
rect 96616 22272 96680 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 81016 21788 81080 21792
rect 81016 21732 81020 21788
rect 81020 21732 81076 21788
rect 81076 21732 81080 21788
rect 81016 21728 81080 21732
rect 81096 21788 81160 21792
rect 81096 21732 81100 21788
rect 81100 21732 81156 21788
rect 81156 21732 81160 21788
rect 81096 21728 81160 21732
rect 81176 21788 81240 21792
rect 81176 21732 81180 21788
rect 81180 21732 81236 21788
rect 81236 21732 81240 21788
rect 81176 21728 81240 21732
rect 81256 21788 81320 21792
rect 81256 21732 81260 21788
rect 81260 21732 81316 21788
rect 81316 21732 81320 21788
rect 81256 21728 81320 21732
rect 111736 21788 111800 21792
rect 111736 21732 111740 21788
rect 111740 21732 111796 21788
rect 111796 21732 111800 21788
rect 111736 21728 111800 21732
rect 111816 21788 111880 21792
rect 111816 21732 111820 21788
rect 111820 21732 111876 21788
rect 111876 21732 111880 21788
rect 111816 21728 111880 21732
rect 111896 21788 111960 21792
rect 111896 21732 111900 21788
rect 111900 21732 111956 21788
rect 111956 21732 111960 21788
rect 111896 21728 111960 21732
rect 111976 21788 112040 21792
rect 111976 21732 111980 21788
rect 111980 21732 112036 21788
rect 112036 21732 112040 21788
rect 111976 21728 112040 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 96376 21244 96440 21248
rect 96376 21188 96380 21244
rect 96380 21188 96436 21244
rect 96436 21188 96440 21244
rect 96376 21184 96440 21188
rect 96456 21244 96520 21248
rect 96456 21188 96460 21244
rect 96460 21188 96516 21244
rect 96516 21188 96520 21244
rect 96456 21184 96520 21188
rect 96536 21244 96600 21248
rect 96536 21188 96540 21244
rect 96540 21188 96596 21244
rect 96596 21188 96600 21244
rect 96536 21184 96600 21188
rect 96616 21244 96680 21248
rect 96616 21188 96620 21244
rect 96620 21188 96676 21244
rect 96676 21188 96680 21244
rect 96616 21184 96680 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 81016 20700 81080 20704
rect 81016 20644 81020 20700
rect 81020 20644 81076 20700
rect 81076 20644 81080 20700
rect 81016 20640 81080 20644
rect 81096 20700 81160 20704
rect 81096 20644 81100 20700
rect 81100 20644 81156 20700
rect 81156 20644 81160 20700
rect 81096 20640 81160 20644
rect 81176 20700 81240 20704
rect 81176 20644 81180 20700
rect 81180 20644 81236 20700
rect 81236 20644 81240 20700
rect 81176 20640 81240 20644
rect 81256 20700 81320 20704
rect 81256 20644 81260 20700
rect 81260 20644 81316 20700
rect 81316 20644 81320 20700
rect 81256 20640 81320 20644
rect 111736 20700 111800 20704
rect 111736 20644 111740 20700
rect 111740 20644 111796 20700
rect 111796 20644 111800 20700
rect 111736 20640 111800 20644
rect 111816 20700 111880 20704
rect 111816 20644 111820 20700
rect 111820 20644 111876 20700
rect 111876 20644 111880 20700
rect 111816 20640 111880 20644
rect 111896 20700 111960 20704
rect 111896 20644 111900 20700
rect 111900 20644 111956 20700
rect 111956 20644 111960 20700
rect 111896 20640 111960 20644
rect 111976 20700 112040 20704
rect 111976 20644 111980 20700
rect 111980 20644 112036 20700
rect 112036 20644 112040 20700
rect 111976 20640 112040 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 96376 20156 96440 20160
rect 96376 20100 96380 20156
rect 96380 20100 96436 20156
rect 96436 20100 96440 20156
rect 96376 20096 96440 20100
rect 96456 20156 96520 20160
rect 96456 20100 96460 20156
rect 96460 20100 96516 20156
rect 96516 20100 96520 20156
rect 96456 20096 96520 20100
rect 96536 20156 96600 20160
rect 96536 20100 96540 20156
rect 96540 20100 96596 20156
rect 96596 20100 96600 20156
rect 96536 20096 96600 20100
rect 96616 20156 96680 20160
rect 96616 20100 96620 20156
rect 96620 20100 96676 20156
rect 96676 20100 96680 20156
rect 96616 20096 96680 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 81016 19612 81080 19616
rect 81016 19556 81020 19612
rect 81020 19556 81076 19612
rect 81076 19556 81080 19612
rect 81016 19552 81080 19556
rect 81096 19612 81160 19616
rect 81096 19556 81100 19612
rect 81100 19556 81156 19612
rect 81156 19556 81160 19612
rect 81096 19552 81160 19556
rect 81176 19612 81240 19616
rect 81176 19556 81180 19612
rect 81180 19556 81236 19612
rect 81236 19556 81240 19612
rect 81176 19552 81240 19556
rect 81256 19612 81320 19616
rect 81256 19556 81260 19612
rect 81260 19556 81316 19612
rect 81316 19556 81320 19612
rect 81256 19552 81320 19556
rect 111736 19612 111800 19616
rect 111736 19556 111740 19612
rect 111740 19556 111796 19612
rect 111796 19556 111800 19612
rect 111736 19552 111800 19556
rect 111816 19612 111880 19616
rect 111816 19556 111820 19612
rect 111820 19556 111876 19612
rect 111876 19556 111880 19612
rect 111816 19552 111880 19556
rect 111896 19612 111960 19616
rect 111896 19556 111900 19612
rect 111900 19556 111956 19612
rect 111956 19556 111960 19612
rect 111896 19552 111960 19556
rect 111976 19612 112040 19616
rect 111976 19556 111980 19612
rect 111980 19556 112036 19612
rect 112036 19556 112040 19612
rect 111976 19552 112040 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 96376 19068 96440 19072
rect 96376 19012 96380 19068
rect 96380 19012 96436 19068
rect 96436 19012 96440 19068
rect 96376 19008 96440 19012
rect 96456 19068 96520 19072
rect 96456 19012 96460 19068
rect 96460 19012 96516 19068
rect 96516 19012 96520 19068
rect 96456 19008 96520 19012
rect 96536 19068 96600 19072
rect 96536 19012 96540 19068
rect 96540 19012 96596 19068
rect 96596 19012 96600 19068
rect 96536 19008 96600 19012
rect 96616 19068 96680 19072
rect 96616 19012 96620 19068
rect 96620 19012 96676 19068
rect 96676 19012 96680 19068
rect 96616 19008 96680 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 81016 18524 81080 18528
rect 81016 18468 81020 18524
rect 81020 18468 81076 18524
rect 81076 18468 81080 18524
rect 81016 18464 81080 18468
rect 81096 18524 81160 18528
rect 81096 18468 81100 18524
rect 81100 18468 81156 18524
rect 81156 18468 81160 18524
rect 81096 18464 81160 18468
rect 81176 18524 81240 18528
rect 81176 18468 81180 18524
rect 81180 18468 81236 18524
rect 81236 18468 81240 18524
rect 81176 18464 81240 18468
rect 81256 18524 81320 18528
rect 81256 18468 81260 18524
rect 81260 18468 81316 18524
rect 81316 18468 81320 18524
rect 81256 18464 81320 18468
rect 111736 18524 111800 18528
rect 111736 18468 111740 18524
rect 111740 18468 111796 18524
rect 111796 18468 111800 18524
rect 111736 18464 111800 18468
rect 111816 18524 111880 18528
rect 111816 18468 111820 18524
rect 111820 18468 111876 18524
rect 111876 18468 111880 18524
rect 111816 18464 111880 18468
rect 111896 18524 111960 18528
rect 111896 18468 111900 18524
rect 111900 18468 111956 18524
rect 111956 18468 111960 18524
rect 111896 18464 111960 18468
rect 111976 18524 112040 18528
rect 111976 18468 111980 18524
rect 111980 18468 112036 18524
rect 112036 18468 112040 18524
rect 111976 18464 112040 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 96376 17980 96440 17984
rect 96376 17924 96380 17980
rect 96380 17924 96436 17980
rect 96436 17924 96440 17980
rect 96376 17920 96440 17924
rect 96456 17980 96520 17984
rect 96456 17924 96460 17980
rect 96460 17924 96516 17980
rect 96516 17924 96520 17980
rect 96456 17920 96520 17924
rect 96536 17980 96600 17984
rect 96536 17924 96540 17980
rect 96540 17924 96596 17980
rect 96596 17924 96600 17980
rect 96536 17920 96600 17924
rect 96616 17980 96680 17984
rect 96616 17924 96620 17980
rect 96620 17924 96676 17980
rect 96676 17924 96680 17980
rect 96616 17920 96680 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 81016 17436 81080 17440
rect 81016 17380 81020 17436
rect 81020 17380 81076 17436
rect 81076 17380 81080 17436
rect 81016 17376 81080 17380
rect 81096 17436 81160 17440
rect 81096 17380 81100 17436
rect 81100 17380 81156 17436
rect 81156 17380 81160 17436
rect 81096 17376 81160 17380
rect 81176 17436 81240 17440
rect 81176 17380 81180 17436
rect 81180 17380 81236 17436
rect 81236 17380 81240 17436
rect 81176 17376 81240 17380
rect 81256 17436 81320 17440
rect 81256 17380 81260 17436
rect 81260 17380 81316 17436
rect 81316 17380 81320 17436
rect 81256 17376 81320 17380
rect 111736 17436 111800 17440
rect 111736 17380 111740 17436
rect 111740 17380 111796 17436
rect 111796 17380 111800 17436
rect 111736 17376 111800 17380
rect 111816 17436 111880 17440
rect 111816 17380 111820 17436
rect 111820 17380 111876 17436
rect 111876 17380 111880 17436
rect 111816 17376 111880 17380
rect 111896 17436 111960 17440
rect 111896 17380 111900 17436
rect 111900 17380 111956 17436
rect 111956 17380 111960 17436
rect 111896 17376 111960 17380
rect 111976 17436 112040 17440
rect 111976 17380 111980 17436
rect 111980 17380 112036 17436
rect 112036 17380 112040 17436
rect 111976 17376 112040 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 96376 16892 96440 16896
rect 96376 16836 96380 16892
rect 96380 16836 96436 16892
rect 96436 16836 96440 16892
rect 96376 16832 96440 16836
rect 96456 16892 96520 16896
rect 96456 16836 96460 16892
rect 96460 16836 96516 16892
rect 96516 16836 96520 16892
rect 96456 16832 96520 16836
rect 96536 16892 96600 16896
rect 96536 16836 96540 16892
rect 96540 16836 96596 16892
rect 96596 16836 96600 16892
rect 96536 16832 96600 16836
rect 96616 16892 96680 16896
rect 96616 16836 96620 16892
rect 96620 16836 96676 16892
rect 96676 16836 96680 16892
rect 96616 16832 96680 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 81016 16348 81080 16352
rect 81016 16292 81020 16348
rect 81020 16292 81076 16348
rect 81076 16292 81080 16348
rect 81016 16288 81080 16292
rect 81096 16348 81160 16352
rect 81096 16292 81100 16348
rect 81100 16292 81156 16348
rect 81156 16292 81160 16348
rect 81096 16288 81160 16292
rect 81176 16348 81240 16352
rect 81176 16292 81180 16348
rect 81180 16292 81236 16348
rect 81236 16292 81240 16348
rect 81176 16288 81240 16292
rect 81256 16348 81320 16352
rect 81256 16292 81260 16348
rect 81260 16292 81316 16348
rect 81316 16292 81320 16348
rect 81256 16288 81320 16292
rect 111736 16348 111800 16352
rect 111736 16292 111740 16348
rect 111740 16292 111796 16348
rect 111796 16292 111800 16348
rect 111736 16288 111800 16292
rect 111816 16348 111880 16352
rect 111816 16292 111820 16348
rect 111820 16292 111876 16348
rect 111876 16292 111880 16348
rect 111816 16288 111880 16292
rect 111896 16348 111960 16352
rect 111896 16292 111900 16348
rect 111900 16292 111956 16348
rect 111956 16292 111960 16348
rect 111896 16288 111960 16292
rect 111976 16348 112040 16352
rect 111976 16292 111980 16348
rect 111980 16292 112036 16348
rect 112036 16292 112040 16348
rect 111976 16288 112040 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 96376 15804 96440 15808
rect 96376 15748 96380 15804
rect 96380 15748 96436 15804
rect 96436 15748 96440 15804
rect 96376 15744 96440 15748
rect 96456 15804 96520 15808
rect 96456 15748 96460 15804
rect 96460 15748 96516 15804
rect 96516 15748 96520 15804
rect 96456 15744 96520 15748
rect 96536 15804 96600 15808
rect 96536 15748 96540 15804
rect 96540 15748 96596 15804
rect 96596 15748 96600 15804
rect 96536 15744 96600 15748
rect 96616 15804 96680 15808
rect 96616 15748 96620 15804
rect 96620 15748 96676 15804
rect 96676 15748 96680 15804
rect 96616 15744 96680 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 81016 15260 81080 15264
rect 81016 15204 81020 15260
rect 81020 15204 81076 15260
rect 81076 15204 81080 15260
rect 81016 15200 81080 15204
rect 81096 15260 81160 15264
rect 81096 15204 81100 15260
rect 81100 15204 81156 15260
rect 81156 15204 81160 15260
rect 81096 15200 81160 15204
rect 81176 15260 81240 15264
rect 81176 15204 81180 15260
rect 81180 15204 81236 15260
rect 81236 15204 81240 15260
rect 81176 15200 81240 15204
rect 81256 15260 81320 15264
rect 81256 15204 81260 15260
rect 81260 15204 81316 15260
rect 81316 15204 81320 15260
rect 81256 15200 81320 15204
rect 111736 15260 111800 15264
rect 111736 15204 111740 15260
rect 111740 15204 111796 15260
rect 111796 15204 111800 15260
rect 111736 15200 111800 15204
rect 111816 15260 111880 15264
rect 111816 15204 111820 15260
rect 111820 15204 111876 15260
rect 111876 15204 111880 15260
rect 111816 15200 111880 15204
rect 111896 15260 111960 15264
rect 111896 15204 111900 15260
rect 111900 15204 111956 15260
rect 111956 15204 111960 15260
rect 111896 15200 111960 15204
rect 111976 15260 112040 15264
rect 111976 15204 111980 15260
rect 111980 15204 112036 15260
rect 112036 15204 112040 15260
rect 111976 15200 112040 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 96376 14716 96440 14720
rect 96376 14660 96380 14716
rect 96380 14660 96436 14716
rect 96436 14660 96440 14716
rect 96376 14656 96440 14660
rect 96456 14716 96520 14720
rect 96456 14660 96460 14716
rect 96460 14660 96516 14716
rect 96516 14660 96520 14716
rect 96456 14656 96520 14660
rect 96536 14716 96600 14720
rect 96536 14660 96540 14716
rect 96540 14660 96596 14716
rect 96596 14660 96600 14716
rect 96536 14656 96600 14660
rect 96616 14716 96680 14720
rect 96616 14660 96620 14716
rect 96620 14660 96676 14716
rect 96676 14660 96680 14716
rect 96616 14656 96680 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 81016 14172 81080 14176
rect 81016 14116 81020 14172
rect 81020 14116 81076 14172
rect 81076 14116 81080 14172
rect 81016 14112 81080 14116
rect 81096 14172 81160 14176
rect 81096 14116 81100 14172
rect 81100 14116 81156 14172
rect 81156 14116 81160 14172
rect 81096 14112 81160 14116
rect 81176 14172 81240 14176
rect 81176 14116 81180 14172
rect 81180 14116 81236 14172
rect 81236 14116 81240 14172
rect 81176 14112 81240 14116
rect 81256 14172 81320 14176
rect 81256 14116 81260 14172
rect 81260 14116 81316 14172
rect 81316 14116 81320 14172
rect 81256 14112 81320 14116
rect 111736 14172 111800 14176
rect 111736 14116 111740 14172
rect 111740 14116 111796 14172
rect 111796 14116 111800 14172
rect 111736 14112 111800 14116
rect 111816 14172 111880 14176
rect 111816 14116 111820 14172
rect 111820 14116 111876 14172
rect 111876 14116 111880 14172
rect 111816 14112 111880 14116
rect 111896 14172 111960 14176
rect 111896 14116 111900 14172
rect 111900 14116 111956 14172
rect 111956 14116 111960 14172
rect 111896 14112 111960 14116
rect 111976 14172 112040 14176
rect 111976 14116 111980 14172
rect 111980 14116 112036 14172
rect 112036 14116 112040 14172
rect 111976 14112 112040 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 96376 13628 96440 13632
rect 96376 13572 96380 13628
rect 96380 13572 96436 13628
rect 96436 13572 96440 13628
rect 96376 13568 96440 13572
rect 96456 13628 96520 13632
rect 96456 13572 96460 13628
rect 96460 13572 96516 13628
rect 96516 13572 96520 13628
rect 96456 13568 96520 13572
rect 96536 13628 96600 13632
rect 96536 13572 96540 13628
rect 96540 13572 96596 13628
rect 96596 13572 96600 13628
rect 96536 13568 96600 13572
rect 96616 13628 96680 13632
rect 96616 13572 96620 13628
rect 96620 13572 96676 13628
rect 96676 13572 96680 13628
rect 96616 13568 96680 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 81016 13084 81080 13088
rect 81016 13028 81020 13084
rect 81020 13028 81076 13084
rect 81076 13028 81080 13084
rect 81016 13024 81080 13028
rect 81096 13084 81160 13088
rect 81096 13028 81100 13084
rect 81100 13028 81156 13084
rect 81156 13028 81160 13084
rect 81096 13024 81160 13028
rect 81176 13084 81240 13088
rect 81176 13028 81180 13084
rect 81180 13028 81236 13084
rect 81236 13028 81240 13084
rect 81176 13024 81240 13028
rect 81256 13084 81320 13088
rect 81256 13028 81260 13084
rect 81260 13028 81316 13084
rect 81316 13028 81320 13084
rect 81256 13024 81320 13028
rect 111736 13084 111800 13088
rect 111736 13028 111740 13084
rect 111740 13028 111796 13084
rect 111796 13028 111800 13084
rect 111736 13024 111800 13028
rect 111816 13084 111880 13088
rect 111816 13028 111820 13084
rect 111820 13028 111876 13084
rect 111876 13028 111880 13084
rect 111816 13024 111880 13028
rect 111896 13084 111960 13088
rect 111896 13028 111900 13084
rect 111900 13028 111956 13084
rect 111956 13028 111960 13084
rect 111896 13024 111960 13028
rect 111976 13084 112040 13088
rect 111976 13028 111980 13084
rect 111980 13028 112036 13084
rect 112036 13028 112040 13084
rect 111976 13024 112040 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 96376 12540 96440 12544
rect 96376 12484 96380 12540
rect 96380 12484 96436 12540
rect 96436 12484 96440 12540
rect 96376 12480 96440 12484
rect 96456 12540 96520 12544
rect 96456 12484 96460 12540
rect 96460 12484 96516 12540
rect 96516 12484 96520 12540
rect 96456 12480 96520 12484
rect 96536 12540 96600 12544
rect 96536 12484 96540 12540
rect 96540 12484 96596 12540
rect 96596 12484 96600 12540
rect 96536 12480 96600 12484
rect 96616 12540 96680 12544
rect 96616 12484 96620 12540
rect 96620 12484 96676 12540
rect 96676 12484 96680 12540
rect 96616 12480 96680 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 81016 11996 81080 12000
rect 81016 11940 81020 11996
rect 81020 11940 81076 11996
rect 81076 11940 81080 11996
rect 81016 11936 81080 11940
rect 81096 11996 81160 12000
rect 81096 11940 81100 11996
rect 81100 11940 81156 11996
rect 81156 11940 81160 11996
rect 81096 11936 81160 11940
rect 81176 11996 81240 12000
rect 81176 11940 81180 11996
rect 81180 11940 81236 11996
rect 81236 11940 81240 11996
rect 81176 11936 81240 11940
rect 81256 11996 81320 12000
rect 81256 11940 81260 11996
rect 81260 11940 81316 11996
rect 81316 11940 81320 11996
rect 81256 11936 81320 11940
rect 111736 11996 111800 12000
rect 111736 11940 111740 11996
rect 111740 11940 111796 11996
rect 111796 11940 111800 11996
rect 111736 11936 111800 11940
rect 111816 11996 111880 12000
rect 111816 11940 111820 11996
rect 111820 11940 111876 11996
rect 111876 11940 111880 11996
rect 111816 11936 111880 11940
rect 111896 11996 111960 12000
rect 111896 11940 111900 11996
rect 111900 11940 111956 11996
rect 111956 11940 111960 11996
rect 111896 11936 111960 11940
rect 111976 11996 112040 12000
rect 111976 11940 111980 11996
rect 111980 11940 112036 11996
rect 112036 11940 112040 11996
rect 111976 11936 112040 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 96376 11452 96440 11456
rect 96376 11396 96380 11452
rect 96380 11396 96436 11452
rect 96436 11396 96440 11452
rect 96376 11392 96440 11396
rect 96456 11452 96520 11456
rect 96456 11396 96460 11452
rect 96460 11396 96516 11452
rect 96516 11396 96520 11452
rect 96456 11392 96520 11396
rect 96536 11452 96600 11456
rect 96536 11396 96540 11452
rect 96540 11396 96596 11452
rect 96596 11396 96600 11452
rect 96536 11392 96600 11396
rect 96616 11452 96680 11456
rect 96616 11396 96620 11452
rect 96620 11396 96676 11452
rect 96676 11396 96680 11452
rect 96616 11392 96680 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 81016 10908 81080 10912
rect 81016 10852 81020 10908
rect 81020 10852 81076 10908
rect 81076 10852 81080 10908
rect 81016 10848 81080 10852
rect 81096 10908 81160 10912
rect 81096 10852 81100 10908
rect 81100 10852 81156 10908
rect 81156 10852 81160 10908
rect 81096 10848 81160 10852
rect 81176 10908 81240 10912
rect 81176 10852 81180 10908
rect 81180 10852 81236 10908
rect 81236 10852 81240 10908
rect 81176 10848 81240 10852
rect 81256 10908 81320 10912
rect 81256 10852 81260 10908
rect 81260 10852 81316 10908
rect 81316 10852 81320 10908
rect 81256 10848 81320 10852
rect 111736 10908 111800 10912
rect 111736 10852 111740 10908
rect 111740 10852 111796 10908
rect 111796 10852 111800 10908
rect 111736 10848 111800 10852
rect 111816 10908 111880 10912
rect 111816 10852 111820 10908
rect 111820 10852 111876 10908
rect 111876 10852 111880 10908
rect 111816 10848 111880 10852
rect 111896 10908 111960 10912
rect 111896 10852 111900 10908
rect 111900 10852 111956 10908
rect 111956 10852 111960 10908
rect 111896 10848 111960 10852
rect 111976 10908 112040 10912
rect 111976 10852 111980 10908
rect 111980 10852 112036 10908
rect 112036 10852 112040 10908
rect 111976 10848 112040 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 96376 10364 96440 10368
rect 96376 10308 96380 10364
rect 96380 10308 96436 10364
rect 96436 10308 96440 10364
rect 96376 10304 96440 10308
rect 96456 10364 96520 10368
rect 96456 10308 96460 10364
rect 96460 10308 96516 10364
rect 96516 10308 96520 10364
rect 96456 10304 96520 10308
rect 96536 10364 96600 10368
rect 96536 10308 96540 10364
rect 96540 10308 96596 10364
rect 96596 10308 96600 10364
rect 96536 10304 96600 10308
rect 96616 10364 96680 10368
rect 96616 10308 96620 10364
rect 96620 10308 96676 10364
rect 96676 10308 96680 10364
rect 96616 10304 96680 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 81016 9820 81080 9824
rect 81016 9764 81020 9820
rect 81020 9764 81076 9820
rect 81076 9764 81080 9820
rect 81016 9760 81080 9764
rect 81096 9820 81160 9824
rect 81096 9764 81100 9820
rect 81100 9764 81156 9820
rect 81156 9764 81160 9820
rect 81096 9760 81160 9764
rect 81176 9820 81240 9824
rect 81176 9764 81180 9820
rect 81180 9764 81236 9820
rect 81236 9764 81240 9820
rect 81176 9760 81240 9764
rect 81256 9820 81320 9824
rect 81256 9764 81260 9820
rect 81260 9764 81316 9820
rect 81316 9764 81320 9820
rect 81256 9760 81320 9764
rect 111736 9820 111800 9824
rect 111736 9764 111740 9820
rect 111740 9764 111796 9820
rect 111796 9764 111800 9820
rect 111736 9760 111800 9764
rect 111816 9820 111880 9824
rect 111816 9764 111820 9820
rect 111820 9764 111876 9820
rect 111876 9764 111880 9820
rect 111816 9760 111880 9764
rect 111896 9820 111960 9824
rect 111896 9764 111900 9820
rect 111900 9764 111956 9820
rect 111956 9764 111960 9820
rect 111896 9760 111960 9764
rect 111976 9820 112040 9824
rect 111976 9764 111980 9820
rect 111980 9764 112036 9820
rect 112036 9764 112040 9820
rect 111976 9760 112040 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 96376 9276 96440 9280
rect 96376 9220 96380 9276
rect 96380 9220 96436 9276
rect 96436 9220 96440 9276
rect 96376 9216 96440 9220
rect 96456 9276 96520 9280
rect 96456 9220 96460 9276
rect 96460 9220 96516 9276
rect 96516 9220 96520 9276
rect 96456 9216 96520 9220
rect 96536 9276 96600 9280
rect 96536 9220 96540 9276
rect 96540 9220 96596 9276
rect 96596 9220 96600 9276
rect 96536 9216 96600 9220
rect 96616 9276 96680 9280
rect 96616 9220 96620 9276
rect 96620 9220 96676 9276
rect 96676 9220 96680 9276
rect 96616 9216 96680 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 81016 8732 81080 8736
rect 81016 8676 81020 8732
rect 81020 8676 81076 8732
rect 81076 8676 81080 8732
rect 81016 8672 81080 8676
rect 81096 8732 81160 8736
rect 81096 8676 81100 8732
rect 81100 8676 81156 8732
rect 81156 8676 81160 8732
rect 81096 8672 81160 8676
rect 81176 8732 81240 8736
rect 81176 8676 81180 8732
rect 81180 8676 81236 8732
rect 81236 8676 81240 8732
rect 81176 8672 81240 8676
rect 81256 8732 81320 8736
rect 81256 8676 81260 8732
rect 81260 8676 81316 8732
rect 81316 8676 81320 8732
rect 81256 8672 81320 8676
rect 111736 8732 111800 8736
rect 111736 8676 111740 8732
rect 111740 8676 111796 8732
rect 111796 8676 111800 8732
rect 111736 8672 111800 8676
rect 111816 8732 111880 8736
rect 111816 8676 111820 8732
rect 111820 8676 111876 8732
rect 111876 8676 111880 8732
rect 111816 8672 111880 8676
rect 111896 8732 111960 8736
rect 111896 8676 111900 8732
rect 111900 8676 111956 8732
rect 111956 8676 111960 8732
rect 111896 8672 111960 8676
rect 111976 8732 112040 8736
rect 111976 8676 111980 8732
rect 111980 8676 112036 8732
rect 112036 8676 112040 8732
rect 111976 8672 112040 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 96376 8188 96440 8192
rect 96376 8132 96380 8188
rect 96380 8132 96436 8188
rect 96436 8132 96440 8188
rect 96376 8128 96440 8132
rect 96456 8188 96520 8192
rect 96456 8132 96460 8188
rect 96460 8132 96516 8188
rect 96516 8132 96520 8188
rect 96456 8128 96520 8132
rect 96536 8188 96600 8192
rect 96536 8132 96540 8188
rect 96540 8132 96596 8188
rect 96596 8132 96600 8188
rect 96536 8128 96600 8132
rect 96616 8188 96680 8192
rect 96616 8132 96620 8188
rect 96620 8132 96676 8188
rect 96676 8132 96680 8188
rect 96616 8128 96680 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 81016 7644 81080 7648
rect 81016 7588 81020 7644
rect 81020 7588 81076 7644
rect 81076 7588 81080 7644
rect 81016 7584 81080 7588
rect 81096 7644 81160 7648
rect 81096 7588 81100 7644
rect 81100 7588 81156 7644
rect 81156 7588 81160 7644
rect 81096 7584 81160 7588
rect 81176 7644 81240 7648
rect 81176 7588 81180 7644
rect 81180 7588 81236 7644
rect 81236 7588 81240 7644
rect 81176 7584 81240 7588
rect 81256 7644 81320 7648
rect 81256 7588 81260 7644
rect 81260 7588 81316 7644
rect 81316 7588 81320 7644
rect 81256 7584 81320 7588
rect 111736 7644 111800 7648
rect 111736 7588 111740 7644
rect 111740 7588 111796 7644
rect 111796 7588 111800 7644
rect 111736 7584 111800 7588
rect 111816 7644 111880 7648
rect 111816 7588 111820 7644
rect 111820 7588 111876 7644
rect 111876 7588 111880 7644
rect 111816 7584 111880 7588
rect 111896 7644 111960 7648
rect 111896 7588 111900 7644
rect 111900 7588 111956 7644
rect 111956 7588 111960 7644
rect 111896 7584 111960 7588
rect 111976 7644 112040 7648
rect 111976 7588 111980 7644
rect 111980 7588 112036 7644
rect 112036 7588 112040 7644
rect 111976 7584 112040 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 81016 6556 81080 6560
rect 81016 6500 81020 6556
rect 81020 6500 81076 6556
rect 81076 6500 81080 6556
rect 81016 6496 81080 6500
rect 81096 6556 81160 6560
rect 81096 6500 81100 6556
rect 81100 6500 81156 6556
rect 81156 6500 81160 6556
rect 81096 6496 81160 6500
rect 81176 6556 81240 6560
rect 81176 6500 81180 6556
rect 81180 6500 81236 6556
rect 81236 6500 81240 6556
rect 81176 6496 81240 6500
rect 81256 6556 81320 6560
rect 81256 6500 81260 6556
rect 81260 6500 81316 6556
rect 81316 6500 81320 6556
rect 81256 6496 81320 6500
rect 111736 6556 111800 6560
rect 111736 6500 111740 6556
rect 111740 6500 111796 6556
rect 111796 6500 111800 6556
rect 111736 6496 111800 6500
rect 111816 6556 111880 6560
rect 111816 6500 111820 6556
rect 111820 6500 111876 6556
rect 111876 6500 111880 6556
rect 111816 6496 111880 6500
rect 111896 6556 111960 6560
rect 111896 6500 111900 6556
rect 111900 6500 111956 6556
rect 111956 6500 111960 6556
rect 111896 6496 111960 6500
rect 111976 6556 112040 6560
rect 111976 6500 111980 6556
rect 111980 6500 112036 6556
rect 112036 6500 112040 6556
rect 111976 6496 112040 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 81016 5468 81080 5472
rect 81016 5412 81020 5468
rect 81020 5412 81076 5468
rect 81076 5412 81080 5468
rect 81016 5408 81080 5412
rect 81096 5468 81160 5472
rect 81096 5412 81100 5468
rect 81100 5412 81156 5468
rect 81156 5412 81160 5468
rect 81096 5408 81160 5412
rect 81176 5468 81240 5472
rect 81176 5412 81180 5468
rect 81180 5412 81236 5468
rect 81236 5412 81240 5468
rect 81176 5408 81240 5412
rect 81256 5468 81320 5472
rect 81256 5412 81260 5468
rect 81260 5412 81316 5468
rect 81316 5412 81320 5468
rect 81256 5408 81320 5412
rect 111736 5468 111800 5472
rect 111736 5412 111740 5468
rect 111740 5412 111796 5468
rect 111796 5412 111800 5468
rect 111736 5408 111800 5412
rect 111816 5468 111880 5472
rect 111816 5412 111820 5468
rect 111820 5412 111876 5468
rect 111876 5412 111880 5468
rect 111816 5408 111880 5412
rect 111896 5468 111960 5472
rect 111896 5412 111900 5468
rect 111900 5412 111956 5468
rect 111956 5412 111960 5468
rect 111896 5408 111960 5412
rect 111976 5468 112040 5472
rect 111976 5412 111980 5468
rect 111980 5412 112036 5468
rect 112036 5412 112040 5468
rect 111976 5408 112040 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 81016 4380 81080 4384
rect 81016 4324 81020 4380
rect 81020 4324 81076 4380
rect 81076 4324 81080 4380
rect 81016 4320 81080 4324
rect 81096 4380 81160 4384
rect 81096 4324 81100 4380
rect 81100 4324 81156 4380
rect 81156 4324 81160 4380
rect 81096 4320 81160 4324
rect 81176 4380 81240 4384
rect 81176 4324 81180 4380
rect 81180 4324 81236 4380
rect 81236 4324 81240 4380
rect 81176 4320 81240 4324
rect 81256 4380 81320 4384
rect 81256 4324 81260 4380
rect 81260 4324 81316 4380
rect 81316 4324 81320 4380
rect 81256 4320 81320 4324
rect 111736 4380 111800 4384
rect 111736 4324 111740 4380
rect 111740 4324 111796 4380
rect 111796 4324 111800 4380
rect 111736 4320 111800 4324
rect 111816 4380 111880 4384
rect 111816 4324 111820 4380
rect 111820 4324 111876 4380
rect 111876 4324 111880 4380
rect 111816 4320 111880 4324
rect 111896 4380 111960 4384
rect 111896 4324 111900 4380
rect 111900 4324 111956 4380
rect 111956 4324 111960 4380
rect 111896 4320 111960 4324
rect 111976 4380 112040 4384
rect 111976 4324 111980 4380
rect 111980 4324 112036 4380
rect 112036 4324 112040 4380
rect 111976 4320 112040 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 81016 3292 81080 3296
rect 81016 3236 81020 3292
rect 81020 3236 81076 3292
rect 81076 3236 81080 3292
rect 81016 3232 81080 3236
rect 81096 3292 81160 3296
rect 81096 3236 81100 3292
rect 81100 3236 81156 3292
rect 81156 3236 81160 3292
rect 81096 3232 81160 3236
rect 81176 3292 81240 3296
rect 81176 3236 81180 3292
rect 81180 3236 81236 3292
rect 81236 3236 81240 3292
rect 81176 3232 81240 3236
rect 81256 3292 81320 3296
rect 81256 3236 81260 3292
rect 81260 3236 81316 3292
rect 81316 3236 81320 3292
rect 81256 3232 81320 3236
rect 111736 3292 111800 3296
rect 111736 3236 111740 3292
rect 111740 3236 111796 3292
rect 111796 3236 111800 3292
rect 111736 3232 111800 3236
rect 111816 3292 111880 3296
rect 111816 3236 111820 3292
rect 111820 3236 111876 3292
rect 111876 3236 111880 3292
rect 111816 3232 111880 3236
rect 111896 3292 111960 3296
rect 111896 3236 111900 3292
rect 111900 3236 111956 3292
rect 111956 3236 111960 3292
rect 111896 3232 111960 3236
rect 111976 3292 112040 3296
rect 111976 3236 111980 3292
rect 111980 3236 112036 3292
rect 112036 3236 112040 3292
rect 111976 3232 112040 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 81016 2204 81080 2208
rect 81016 2148 81020 2204
rect 81020 2148 81076 2204
rect 81076 2148 81080 2204
rect 81016 2144 81080 2148
rect 81096 2204 81160 2208
rect 81096 2148 81100 2204
rect 81100 2148 81156 2204
rect 81156 2148 81160 2204
rect 81096 2144 81160 2148
rect 81176 2204 81240 2208
rect 81176 2148 81180 2204
rect 81180 2148 81236 2204
rect 81236 2148 81240 2204
rect 81176 2144 81240 2148
rect 81256 2204 81320 2208
rect 81256 2148 81260 2204
rect 81260 2148 81316 2204
rect 81316 2148 81320 2204
rect 81256 2144 81320 2148
rect 111736 2204 111800 2208
rect 111736 2148 111740 2204
rect 111740 2148 111796 2204
rect 111796 2148 111800 2204
rect 111736 2144 111800 2148
rect 111816 2204 111880 2208
rect 111816 2148 111820 2204
rect 111820 2148 111876 2204
rect 111876 2148 111880 2204
rect 111816 2144 111880 2148
rect 111896 2204 111960 2208
rect 111896 2148 111900 2204
rect 111900 2148 111956 2204
rect 111956 2148 111960 2204
rect 111896 2144 111960 2148
rect 111976 2204 112040 2208
rect 111976 2148 111980 2204
rect 111980 2148 112036 2204
rect 112036 2148 112040 2204
rect 111976 2144 112040 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 37024 50608 37584
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 37568 65968 37584
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
rect 81008 37024 81328 37584
rect 81008 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81328 37024
rect 81008 35936 81328 36960
rect 81008 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81328 35936
rect 81008 34848 81328 35872
rect 81008 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81328 34848
rect 81008 33760 81328 34784
rect 81008 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81328 33760
rect 81008 32672 81328 33696
rect 81008 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81328 32672
rect 81008 31584 81328 32608
rect 81008 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81328 31584
rect 81008 30496 81328 31520
rect 81008 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81328 30496
rect 81008 29408 81328 30432
rect 81008 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81328 29408
rect 81008 28320 81328 29344
rect 81008 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81328 28320
rect 81008 27232 81328 28256
rect 81008 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81328 27232
rect 81008 26144 81328 27168
rect 81008 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81328 26144
rect 81008 25056 81328 26080
rect 81008 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81328 25056
rect 81008 23968 81328 24992
rect 81008 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81328 23968
rect 81008 22880 81328 23904
rect 81008 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81328 22880
rect 81008 21792 81328 22816
rect 81008 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81328 21792
rect 81008 20704 81328 21728
rect 81008 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81328 20704
rect 81008 19616 81328 20640
rect 81008 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81328 19616
rect 81008 18528 81328 19552
rect 81008 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81328 18528
rect 81008 17440 81328 18464
rect 81008 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81328 17440
rect 81008 16352 81328 17376
rect 81008 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81328 16352
rect 81008 15264 81328 16288
rect 81008 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81328 15264
rect 81008 14176 81328 15200
rect 81008 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81328 14176
rect 81008 13088 81328 14112
rect 81008 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81328 13088
rect 81008 12000 81328 13024
rect 81008 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81328 12000
rect 81008 10912 81328 11936
rect 81008 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81328 10912
rect 81008 9824 81328 10848
rect 81008 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81328 9824
rect 81008 8736 81328 9760
rect 81008 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81328 8736
rect 81008 7648 81328 8672
rect 81008 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81328 7648
rect 81008 6560 81328 7584
rect 81008 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81328 6560
rect 81008 5472 81328 6496
rect 81008 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81328 5472
rect 81008 4384 81328 5408
rect 81008 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81328 4384
rect 81008 3296 81328 4320
rect 81008 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81328 3296
rect 81008 2208 81328 3232
rect 81008 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81328 2208
rect 81008 2128 81328 2144
rect 96368 37568 96688 37584
rect 96368 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96688 37568
rect 96368 36480 96688 37504
rect 96368 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96688 36480
rect 96368 35392 96688 36416
rect 96368 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96688 35392
rect 96368 34304 96688 35328
rect 96368 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96688 34304
rect 96368 33216 96688 34240
rect 96368 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96688 33216
rect 96368 32128 96688 33152
rect 96368 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96688 32128
rect 96368 31040 96688 32064
rect 96368 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96688 31040
rect 96368 29952 96688 30976
rect 96368 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96688 29952
rect 96368 28864 96688 29888
rect 96368 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96688 28864
rect 96368 27776 96688 28800
rect 96368 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96688 27776
rect 96368 26688 96688 27712
rect 96368 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96688 26688
rect 96368 25600 96688 26624
rect 96368 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96688 25600
rect 96368 24512 96688 25536
rect 96368 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96688 24512
rect 96368 23424 96688 24448
rect 96368 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96688 23424
rect 96368 22336 96688 23360
rect 96368 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96688 22336
rect 96368 21248 96688 22272
rect 96368 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96688 21248
rect 96368 20160 96688 21184
rect 96368 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96688 20160
rect 96368 19072 96688 20096
rect 96368 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96688 19072
rect 96368 17984 96688 19008
rect 96368 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96688 17984
rect 96368 16896 96688 17920
rect 96368 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96688 16896
rect 96368 15808 96688 16832
rect 96368 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96688 15808
rect 96368 14720 96688 15744
rect 96368 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96688 14720
rect 96368 13632 96688 14656
rect 96368 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96688 13632
rect 96368 12544 96688 13568
rect 96368 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96688 12544
rect 96368 11456 96688 12480
rect 96368 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96688 11456
rect 96368 10368 96688 11392
rect 96368 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96688 10368
rect 96368 9280 96688 10304
rect 96368 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96688 9280
rect 96368 8192 96688 9216
rect 96368 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96688 8192
rect 96368 7104 96688 8128
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 4928 96688 5952
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 111728 37024 112048 37584
rect 111728 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112048 37024
rect 111728 35936 112048 36960
rect 111728 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112048 35936
rect 111728 34848 112048 35872
rect 111728 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112048 34848
rect 111728 33760 112048 34784
rect 111728 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112048 33760
rect 111728 32672 112048 33696
rect 111728 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112048 32672
rect 111728 31584 112048 32608
rect 111728 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112048 31584
rect 111728 30496 112048 31520
rect 111728 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112048 30496
rect 111728 29408 112048 30432
rect 111728 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112048 29408
rect 111728 28320 112048 29344
rect 111728 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112048 28320
rect 111728 27232 112048 28256
rect 111728 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112048 27232
rect 111728 26144 112048 27168
rect 111728 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112048 26144
rect 111728 25056 112048 26080
rect 111728 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112048 25056
rect 111728 23968 112048 24992
rect 111728 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112048 23968
rect 111728 22880 112048 23904
rect 111728 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112048 22880
rect 111728 21792 112048 22816
rect 111728 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112048 21792
rect 111728 20704 112048 21728
rect 111728 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112048 20704
rect 111728 19616 112048 20640
rect 111728 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112048 19616
rect 111728 18528 112048 19552
rect 111728 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112048 18528
rect 111728 17440 112048 18464
rect 111728 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112048 17440
rect 111728 16352 112048 17376
rect 111728 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112048 16352
rect 111728 15264 112048 16288
rect 111728 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112048 15264
rect 111728 14176 112048 15200
rect 111728 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112048 14176
rect 111728 13088 112048 14112
rect 111728 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112048 13088
rect 111728 12000 112048 13024
rect 111728 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112048 12000
rect 111728 10912 112048 11936
rect 111728 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112048 10912
rect 111728 9824 112048 10848
rect 111728 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112048 9824
rect 111728 8736 112048 9760
rect 111728 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112048 8736
rect 111728 7648 112048 8672
rect 111728 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112048 7648
rect 111728 6560 112048 7584
rect 111728 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112048 6560
rect 111728 5472 112048 6496
rect 111728 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112048 5472
rect 111728 4384 112048 5408
rect 111728 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112048 4384
rect 111728 3296 112048 4320
rect 111728 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112048 3296
rect 111728 2208 112048 3232
rect 111728 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112048 2208
rect 111728 2128 112048 2144
use sky130_fd_sc_hd__decap_8  FILLER_0_19 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1644511149
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60
timestamp 1644511149
transform 1 0 6624 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_116
timestamp 1644511149
transform 1 0 11776 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_122
timestamp 1644511149
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1644511149
transform 1 0 13524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1644511149
transform 1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_213
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_232
timestamp 1644511149
transform 1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_239
timestamp 1644511149
transform 1 0 23092 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1644511149
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_291
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_302
timestamp 1644511149
transform 1 0 28888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1644511149
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_315
timestamp 1644511149
transform 1 0 30084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_319
timestamp 1644511149
transform 1 0 30452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1644511149
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_330
timestamp 1644511149
transform 1 0 31464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_343
timestamp 1644511149
transform 1 0 32660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1644511149
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1644511149
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_380
timestamp 1644511149
transform 1 0 36064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_397
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1644511149
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_408
timestamp 1644511149
transform 1 0 38640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_425
timestamp 1644511149
transform 1 0 40204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_428
timestamp 1644511149
transform 1 0 40480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_434
timestamp 1644511149
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_441
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1644511149
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_464
timestamp 1644511149
transform 1 0 43792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1644511149
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1644511149
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_482
timestamp 1644511149
transform 1 0 45448 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_491
timestamp 1644511149
transform 1 0 46276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_510
timestamp 1644511149
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1644511149
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_543
timestamp 1644511149
transform 1 0 51060 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_551
timestamp 1644511149
transform 1 0 51796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_556
timestamp 1644511149
transform 1 0 52256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_566
timestamp 1644511149
transform 1 0 53176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1644511149
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1644511149
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1644511149
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_621
timestamp 1644511149
transform 1 0 58236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_633
timestamp 1644511149
transform 1 0 59340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_640
timestamp 1644511149
transform 1 0 59984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_648
timestamp 1644511149
transform 1 0 60720 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_656
timestamp 1644511149
transform 1 0 61456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_662
timestamp 1644511149
transform 1 0 62008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_670
timestamp 1644511149
transform 1 0 62744 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_678
timestamp 1644511149
transform 1 0 63480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_685
timestamp 1644511149
transform 1 0 64124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_692
timestamp 1644511149
transform 1 0 64768 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_706
timestamp 1644511149
transform 1 0 66056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_715
timestamp 1644511149
transform 1 0 66884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_722
timestamp 1644511149
transform 1 0 67528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_729
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_737
timestamp 1644511149
transform 1 0 68908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_744
timestamp 1644511149
transform 1 0 69552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_751
timestamp 1644511149
transform 1 0 70196 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 1644511149
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_760
timestamp 1644511149
transform 1 0 71024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_769
timestamp 1644511149
transform 1 0 71852 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_778
timestamp 1644511149
transform 1 0 72680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_790
timestamp 1644511149
transform 1 0 73784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_803
timestamp 1644511149
transform 1 0 74980 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 1644511149
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_817
timestamp 1644511149
transform 1 0 76268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_830
timestamp 1644511149
transform 1 0 77464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_838
timestamp 1644511149
transform 1 0 78200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_845
timestamp 1644511149
transform 1 0 78844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_852
timestamp 1644511149
transform 1 0 79488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_859
timestamp 1644511149
transform 1 0 80132 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_867
timestamp 1644511149
transform 1 0 80868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_869
timestamp 1644511149
transform 1 0 81052 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_874
timestamp 1644511149
transform 1 0 81512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_883
timestamp 1644511149
transform 1 0 82340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_892
timestamp 1644511149
transform 1 0 83168 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_900
timestamp 1644511149
transform 1 0 83904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_904
timestamp 1644511149
transform 1 0 84272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_908
timestamp 1644511149
transform 1 0 84640 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_918
timestamp 1644511149
transform 1 0 85560 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_925
timestamp 1644511149
transform 1 0 86204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_933
timestamp 1644511149
transform 1 0 86940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_941
timestamp 1644511149
transform 1 0 87676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_947
timestamp 1644511149
transform 1 0 88228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_951
timestamp 1644511149
transform 1 0 88596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_956
timestamp 1644511149
transform 1 0 89056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_963
timestamp 1644511149
transform 1 0 89700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_976
timestamp 1644511149
transform 1 0 90896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_986
timestamp 1644511149
transform 1 0 91816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_995
timestamp 1644511149
transform 1 0 92644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1002
timestamp 1644511149
transform 1 0 93288 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1012
timestamp 1644511149
transform 1 0 94208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1019
timestamp 1644511149
transform 1 0 94852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1030
timestamp 1644511149
transform 1 0 95864 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1042
timestamp 1644511149
transform 1 0 96968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1051
timestamp 1644511149
transform 1 0 97796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1058
timestamp 1644511149
transform 1 0 98440 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1081
timestamp 1644511149
transform 1 0 100556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1086
timestamp 1644511149
transform 1 0 101016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1090
timestamp 1644511149
transform 1 0 101384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1097
timestamp 1644511149
transform 1 0 102028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1101
timestamp 1644511149
transform 1 0 102396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1109
timestamp 1644511149
transform 1 0 103132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1113
timestamp 1644511149
transform 1 0 103500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1117
timestamp 1644511149
transform 1 0 103868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1121
timestamp 1644511149
transform 1 0 104236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1141
timestamp 1644511149
transform 1 0 106076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1147
timestamp 1644511149
transform 1 0 106628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1149
timestamp 1644511149
transform 1 0 106812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1161
timestamp 1644511149
transform 1 0 107916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1168
timestamp 1644511149
transform 1 0 108560 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1186
timestamp 1644511149
transform 1 0 110216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1193
timestamp 1644511149
transform 1 0 110860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1208
timestamp 1644511149
transform 1 0 112240 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1216
timestamp 1644511149
transform 1 0 112976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1222
timestamp 1644511149
transform 1 0 113528 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1230
timestamp 1644511149
transform 1 0 114264 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1237
timestamp 1644511149
transform 1 0 114908 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1243
timestamp 1644511149
transform 1 0 115460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1254
timestamp 1644511149
transform 1 0 116472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1265
timestamp 1644511149
transform 1 0 117484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1273
timestamp 1644511149
transform 1 0 118220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1644511149
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_230
timestamp 1644511149
transform 1 0 22264 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_242
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_254
timestamp 1644511149
transform 1 0 24472 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_266
timestamp 1644511149
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1644511149
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_308
timestamp 1644511149
transform 1 0 29440 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_320
timestamp 1644511149
transform 1 0 30544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_328
timestamp 1644511149
transform 1 0 31280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1644511149
transform 1 0 32568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1644511149
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_369
timestamp 1644511149
transform 1 0 35052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1644511149
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_396
timestamp 1644511149
transform 1 0 37536 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_408
timestamp 1644511149
transform 1 0 38640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_416
timestamp 1644511149
transform 1 0 39376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_426
timestamp 1644511149
transform 1 0 40296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1644511149
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1644511149
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_462
timestamp 1644511149
transform 1 0 43608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_469
timestamp 1644511149
transform 1 0 44252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_481
timestamp 1644511149
transform 1 0 45356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_493
timestamp 1644511149
transform 1 0 46460 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_501
timestamp 1644511149
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_510
timestamp 1644511149
transform 1 0 48024 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_522
timestamp 1644511149
transform 1 0 49128 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_530
timestamp 1644511149
transform 1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_539
timestamp 1644511149
transform 1 0 50692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_546
timestamp 1644511149
transform 1 0 51336 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_552
timestamp 1644511149
transform 1 0 51888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_556
timestamp 1644511149
transform 1 0 52256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_568
timestamp 1644511149
transform 1 0 53360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_580
timestamp 1644511149
transform 1 0 54464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_587
timestamp 1644511149
transform 1 0 55108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_593
timestamp 1644511149
transform 1 0 55660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1644511149
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_608
timestamp 1644511149
transform 1 0 57040 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_620
timestamp 1644511149
transform 1 0 58144 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_632
timestamp 1644511149
transform 1 0 59248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_639
timestamp 1644511149
transform 1 0 59892 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_651
timestamp 1644511149
transform 1 0 60996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_663
timestamp 1644511149
transform 1 0 62100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1644511149
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_676
timestamp 1644511149
transform 1 0 63296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_688
timestamp 1644511149
transform 1 0 64400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_696
timestamp 1644511149
transform 1 0 65136 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_700
timestamp 1644511149
transform 1 0 65504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_706
timestamp 1644511149
transform 1 0 66056 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_713
timestamp 1644511149
transform 1 0 66700 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_725
timestamp 1644511149
transform 1 0 67804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_733
timestamp 1644511149
transform 1 0 68540 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_751
timestamp 1644511149
transform 1 0 70196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_761
timestamp 1644511149
transform 1 0 71116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_773
timestamp 1644511149
transform 1 0 72220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_781
timestamp 1644511149
transform 1 0 72956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_785
timestamp 1644511149
transform 1 0 73324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_792
timestamp 1644511149
transform 1 0 73968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_800
timestamp 1644511149
transform 1 0 74704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_807
timestamp 1644511149
transform 1 0 75348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_815
timestamp 1644511149
transform 1 0 76084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_821
timestamp 1644511149
transform 1 0 76636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_830
timestamp 1644511149
transform 1 0 77464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_838
timestamp 1644511149
transform 1 0 78200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_841
timestamp 1644511149
transform 1 0 78476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_853
timestamp 1644511149
transform 1 0 79580 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_864
timestamp 1644511149
transform 1 0 80592 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_876
timestamp 1644511149
transform 1 0 81696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_882
timestamp 1644511149
transform 1 0 82248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_894
timestamp 1644511149
transform 1 0 83352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_903
timestamp 1644511149
transform 1 0 84180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_915
timestamp 1644511149
transform 1 0 85284 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_926
timestamp 1644511149
transform 1 0 86296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_930
timestamp 1644511149
transform 1 0 86664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_934
timestamp 1644511149
transform 1 0 87032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_948
timestamp 1644511149
transform 1 0 88320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_953
timestamp 1644511149
transform 1 0 88780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_962
timestamp 1644511149
transform 1 0 89608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_966
timestamp 1644511149
transform 1 0 89976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_973
timestamp 1644511149
transform 1 0 90620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_980
timestamp 1644511149
transform 1 0 91264 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_986
timestamp 1644511149
transform 1 0 91816 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_993
timestamp 1644511149
transform 1 0 92460 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1005
timestamp 1644511149
transform 1 0 93564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1025
timestamp 1644511149
transform 1 0 95404 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1033
timestamp 1644511149
transform 1 0 96140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1039
timestamp 1644511149
transform 1 0 96692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1047
timestamp 1644511149
transform 1 0 97428 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1059
timestamp 1644511149
transform 1 0 98532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1063
timestamp 1644511149
transform 1 0 98900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1065
timestamp 1644511149
transform 1 0 99084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1069
timestamp 1644511149
transform 1 0 99452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1074
timestamp 1644511149
transform 1 0 99912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1078
timestamp 1644511149
transform 1 0 100280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1088
timestamp 1644511149
transform 1 0 101200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1100
timestamp 1644511149
transform 1 0 102304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1112
timestamp 1644511149
transform 1 0 103408 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1125
timestamp 1644511149
transform 1 0 104604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1135
timestamp 1644511149
transform 1 0 105524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1147
timestamp 1644511149
transform 1 0 106628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1153
timestamp 1644511149
transform 1 0 107180 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1170
timestamp 1644511149
transform 1 0 108744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1177
timestamp 1644511149
transform 1 0 109388 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1189
timestamp 1644511149
transform 1 0 110492 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1196
timestamp 1644511149
transform 1 0 111136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1216
timestamp 1644511149
transform 1 0 112976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1223
timestamp 1644511149
transform 1 0 113620 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1644511149
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1233
timestamp 1644511149
transform 1 0 114540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1240
timestamp 1644511149
transform 1 0 115184 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_1252
timestamp 1644511149
transform 1 0 116288 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1264
timestamp 1644511149
transform 1 0 117392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1268
timestamp 1644511149
transform 1 0 117760 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1273
timestamp 1644511149
transform 1 0 118220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_11
timestamp 1644511149
transform 1 0 2116 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1644511149
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1644511149
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1644511149
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_206
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_218
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1644511149
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_395
timestamp 1644511149
transform 1 0 37444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_400
timestamp 1644511149
transform 1 0 37904 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_404
timestamp 1644511149
transform 1 0 38272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1644511149
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1644511149
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1644511149
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_495
timestamp 1644511149
transform 1 0 46644 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_508
timestamp 1644511149
transform 1 0 47840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1644511149
transform 1 0 48944 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_537
timestamp 1644511149
transform 1 0 50508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_549
timestamp 1644511149
transform 1 0 51612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_564
timestamp 1644511149
transform 1 0 52992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1644511149
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_595
timestamp 1644511149
transform 1 0 55844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_602
timestamp 1644511149
transform 1 0 56488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_614
timestamp 1644511149
transform 1 0 57592 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_626
timestamp 1644511149
transform 1 0 58696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_634
timestamp 1644511149
transform 1 0 59432 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_642
timestamp 1644511149
transform 1 0 60168 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_657
timestamp 1644511149
transform 1 0 61548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_667
timestamp 1644511149
transform 1 0 62468 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_679
timestamp 1644511149
transform 1 0 63572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_683
timestamp 1644511149
transform 1 0 63940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_690
timestamp 1644511149
transform 1 0 64584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_698
timestamp 1644511149
transform 1 0 65320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_714
timestamp 1644511149
transform 1 0 66792 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_722
timestamp 1644511149
transform 1 0 67528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_733
timestamp 1644511149
transform 1 0 68540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_745
timestamp 1644511149
transform 1 0 69644 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_753
timestamp 1644511149
transform 1 0 70380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_757
timestamp 1644511149
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_769
timestamp 1644511149
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_781
timestamp 1644511149
transform 1 0 72956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_789
timestamp 1644511149
transform 1 0 73692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_795
timestamp 1644511149
transform 1 0 74244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_807
timestamp 1644511149
transform 1 0 75348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1644511149
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_813
timestamp 1644511149
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_825
timestamp 1644511149
transform 1 0 77004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_837
timestamp 1644511149
transform 1 0 78108 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_849
timestamp 1644511149
transform 1 0 79212 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 1644511149
transform 1 0 80316 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 1644511149
transform 1 0 80868 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_869
timestamp 1644511149
transform 1 0 81052 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_881
timestamp 1644511149
transform 1 0 82156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_893
timestamp 1644511149
transform 1 0 83260 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_901
timestamp 1644511149
transform 1 0 83996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_913
timestamp 1644511149
transform 1 0 85100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_921
timestamp 1644511149
transform 1 0 85836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_941
timestamp 1644511149
transform 1 0 87676 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_949
timestamp 1644511149
transform 1 0 88412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_954
timestamp 1644511149
transform 1 0 88872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_958
timestamp 1644511149
transform 1 0 89240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_962
timestamp 1644511149
transform 1 0 89608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_976
timestamp 1644511149
transform 1 0 90896 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_981
timestamp 1644511149
transform 1 0 91356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_997
timestamp 1644511149
transform 1 0 92828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1016
timestamp 1644511149
transform 1 0 94576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1023
timestamp 1644511149
transform 1 0 95220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1035
timestamp 1644511149
transform 1 0 96324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1037
timestamp 1644511149
transform 1 0 96508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1047
timestamp 1644511149
transform 1 0 97428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1057
timestamp 1644511149
transform 1 0 98348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1067
timestamp 1644511149
transform 1 0 99268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1075
timestamp 1644511149
transform 1 0 100004 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1079
timestamp 1644511149
transform 1 0 100372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1644511149
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1101
timestamp 1644511149
transform 1 0 102396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1113
timestamp 1644511149
transform 1 0 103500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1125
timestamp 1644511149
transform 1 0 104604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1137
timestamp 1644511149
transform 1 0 105708 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1145
timestamp 1644511149
transform 1 0 106444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1149
timestamp 1644511149
transform 1 0 106812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1153
timestamp 1644511149
transform 1 0 107180 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1163
timestamp 1644511149
transform 1 0 108100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1170
timestamp 1644511149
transform 1 0 108744 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1182
timestamp 1644511149
transform 1 0 109848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1194
timestamp 1644511149
transform 1 0 110952 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1202
timestamp 1644511149
transform 1 0 111688 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1214
timestamp 1644511149
transform 1 0 112792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1226
timestamp 1644511149
transform 1 0 113896 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1238
timestamp 1644511149
transform 1 0 115000 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1250
timestamp 1644511149
transform 1 0 116104 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1258
timestamp 1644511149
transform 1 0 116840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1261
timestamp 1644511149
transform 1 0 117116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1273
timestamp 1644511149
transform 1 0 118220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_97
timestamp 1644511149
transform 1 0 10028 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_201
timestamp 1644511149
transform 1 0 19596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_207
timestamp 1644511149
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1644511149
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_233
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_240
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_264
timestamp 1644511149
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_299
timestamp 1644511149
transform 1 0 28612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_423
timestamp 1644511149
transform 1 0 40020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_435
timestamp 1644511149
transform 1 0 41124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_653
timestamp 1644511149
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1644511149
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1644511149
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_678
timestamp 1644511149
transform 1 0 63480 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_690
timestamp 1644511149
transform 1 0 64584 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_702
timestamp 1644511149
transform 1 0 65688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_714
timestamp 1644511149
transform 1 0 66792 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_726
timestamp 1644511149
transform 1 0 67896 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_734
timestamp 1644511149
transform 1 0 68632 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_746
timestamp 1644511149
transform 1 0 69736 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_758
timestamp 1644511149
transform 1 0 70840 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_770
timestamp 1644511149
transform 1 0 71944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_780
timestamp 1644511149
transform 1 0 72864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_785
timestamp 1644511149
transform 1 0 73324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_789
timestamp 1644511149
transform 1 0 73692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_795
timestamp 1644511149
transform 1 0 74244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_807
timestamp 1644511149
transform 1 0 75348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_819
timestamp 1644511149
transform 1 0 76452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_827
timestamp 1644511149
transform 1 0 77188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_834
timestamp 1644511149
transform 1 0 77832 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_841
timestamp 1644511149
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_853
timestamp 1644511149
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_865
timestamp 1644511149
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_877
timestamp 1644511149
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1644511149
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1644511149
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_897
timestamp 1644511149
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_909
timestamp 1644511149
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_921
timestamp 1644511149
transform 1 0 85836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_926
timestamp 1644511149
transform 1 0 86296 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_930
timestamp 1644511149
transform 1 0 86664 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_941
timestamp 1644511149
transform 1 0 87676 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_949
timestamp 1644511149
transform 1 0 88412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_953
timestamp 1644511149
transform 1 0 88780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_960
timestamp 1644511149
transform 1 0 89424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_968
timestamp 1644511149
transform 1 0 90160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_973
timestamp 1644511149
transform 1 0 90620 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_980
timestamp 1644511149
transform 1 0 91264 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_992
timestamp 1644511149
transform 1 0 92368 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1004
timestamp 1644511149
transform 1 0 93472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1018
timestamp 1644511149
transform 1 0 94760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1030
timestamp 1644511149
transform 1 0 95864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1042
timestamp 1644511149
transform 1 0 96968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1051
timestamp 1644511149
transform 1 0 97796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1063
timestamp 1644511149
transform 1 0 98900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1065
timestamp 1644511149
transform 1 0 99084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1073
timestamp 1644511149
transform 1 0 99820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1081
timestamp 1644511149
transform 1 0 100556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1095
timestamp 1644511149
transform 1 0 101844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1107
timestamp 1644511149
transform 1 0 102948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1119
timestamp 1644511149
transform 1 0 104052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1124
timestamp 1644511149
transform 1 0 104512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1131
timestamp 1644511149
transform 1 0 105156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1143
timestamp 1644511149
transform 1 0 106260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1151
timestamp 1644511149
transform 1 0 106996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1168
timestamp 1644511149
transform 1 0 108560 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1177
timestamp 1644511149
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1189
timestamp 1644511149
transform 1 0 110492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1207
timestamp 1644511149
transform 1 0 112148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1219
timestamp 1644511149
transform 1 0 113252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1644511149
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1233
timestamp 1644511149
transform 1 0 114540 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1245
timestamp 1644511149
transform 1 0 115644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1257
timestamp 1644511149
transform 1 0 116748 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1273
timestamp 1644511149
transform 1 0 118220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1644511149
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_108
timestamp 1644511149
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_120
timestamp 1644511149
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_132
timestamp 1644511149
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_235
timestamp 1644511149
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_247
timestamp 1644511149
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_285
timestamp 1644511149
transform 1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1644511149
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1644511149
transform 1 0 29808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1644511149
transform 1 0 30912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_336
timestamp 1644511149
transform 1 0 32016 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_348
timestamp 1644511149
transform 1 0 33120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_521
timestamp 1644511149
transform 1 0 49036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_527
timestamp 1644511149
transform 1 0 49588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_538
timestamp 1644511149
transform 1 0 50600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_550
timestamp 1644511149
transform 1 0 51704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_558
timestamp 1644511149
transform 1 0 52440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_565
timestamp 1644511149
transform 1 0 53084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_577
timestamp 1644511149
transform 1 0 54188 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_585
timestamp 1644511149
transform 1 0 54924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_674
timestamp 1644511149
transform 1 0 63112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_686
timestamp 1644511149
transform 1 0 64216 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_698
timestamp 1644511149
transform 1 0 65320 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_741
timestamp 1644511149
transform 1 0 69276 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_753
timestamp 1644511149
transform 1 0 70380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_757
timestamp 1644511149
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_769
timestamp 1644511149
transform 1 0 71852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_777
timestamp 1644511149
transform 1 0 72588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_794
timestamp 1644511149
transform 1 0 74152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_806
timestamp 1644511149
transform 1 0 75256 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_813
timestamp 1644511149
transform 1 0 75900 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_827
timestamp 1644511149
transform 1 0 77188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_839
timestamp 1644511149
transform 1 0 78292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_851
timestamp 1644511149
transform 1 0 79396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_863
timestamp 1644511149
transform 1 0 80500 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1644511149
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_869
timestamp 1644511149
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_881
timestamp 1644511149
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_893
timestamp 1644511149
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_905
timestamp 1644511149
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1644511149
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1644511149
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_925
timestamp 1644511149
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_937
timestamp 1644511149
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_949
timestamp 1644511149
transform 1 0 88412 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_957
timestamp 1644511149
transform 1 0 89148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_976
timestamp 1644511149
transform 1 0 90896 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_981
timestamp 1644511149
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_993
timestamp 1644511149
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1005
timestamp 1644511149
transform 1 0 93564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1014
timestamp 1644511149
transform 1 0 94392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1026
timestamp 1644511149
transform 1 0 95496 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1034
timestamp 1644511149
transform 1 0 96232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1037
timestamp 1644511149
transform 1 0 96508 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1043
timestamp 1644511149
transform 1 0 97060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1050
timestamp 1644511149
transform 1 0 97704 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1062
timestamp 1644511149
transform 1 0 98808 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_1074
timestamp 1644511149
transform 1 0 99912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1080
timestamp 1644511149
transform 1 0 100464 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1093
timestamp 1644511149
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1105
timestamp 1644511149
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1117
timestamp 1644511149
transform 1 0 103868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1123
timestamp 1644511149
transform 1 0 104420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1130
timestamp 1644511149
transform 1 0 105064 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1142
timestamp 1644511149
transform 1 0 106168 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1149
timestamp 1644511149
transform 1 0 106812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1156
timestamp 1644511149
transform 1 0 107456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1168
timestamp 1644511149
transform 1 0 108560 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1180
timestamp 1644511149
transform 1 0 109664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1192
timestamp 1644511149
transform 1 0 110768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1199
timestamp 1644511149
transform 1 0 111412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1644511149
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1214
timestamp 1644511149
transform 1 0 112792 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1226
timestamp 1644511149
transform 1 0 113896 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1238
timestamp 1644511149
transform 1 0 115000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1250
timestamp 1644511149
transform 1 0 116104 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1258
timestamp 1644511149
transform 1 0 116840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1261
timestamp 1644511149
transform 1 0 117116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1273
timestamp 1644511149
transform 1 0 118220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1644511149
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1644511149
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1644511149
transform 1 0 17940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_234
timestamp 1644511149
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_238
timestamp 1644511149
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_250
timestamp 1644511149
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1644511149
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1644511149
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_304
timestamp 1644511149
transform 1 0 29072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_316
timestamp 1644511149
transform 1 0 30176 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1644511149
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_410
timestamp 1644511149
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_423
timestamp 1644511149
transform 1 0 40020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_435
timestamp 1644511149
transform 1 0 41124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_513
timestamp 1644511149
transform 1 0 48300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_532
timestamp 1644511149
transform 1 0 50048 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_545
timestamp 1644511149
transform 1 0 51244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_557
timestamp 1644511149
transform 1 0 52348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_569
timestamp 1644511149
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_576
timestamp 1644511149
transform 1 0 54096 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_588
timestamp 1644511149
transform 1 0 55200 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_600
timestamp 1644511149
transform 1 0 56304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_612
timestamp 1644511149
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_676
timestamp 1644511149
transform 1 0 63296 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_682
timestamp 1644511149
transform 1 0 63848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_692
timestamp 1644511149
transform 1 0 64768 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_704
timestamp 1644511149
transform 1 0 65872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_716
timestamp 1644511149
transform 1 0 66976 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_736
timestamp 1644511149
transform 1 0 68816 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_748
timestamp 1644511149
transform 1 0 69920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_758
timestamp 1644511149
transform 1 0 70840 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_770
timestamp 1644511149
transform 1 0 71944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_782
timestamp 1644511149
transform 1 0 73048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_785
timestamp 1644511149
transform 1 0 73324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_789
timestamp 1644511149
transform 1 0 73692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_801
timestamp 1644511149
transform 1 0 74796 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_807
timestamp 1644511149
transform 1 0 75348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_810
timestamp 1644511149
transform 1 0 75624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_821
timestamp 1644511149
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1644511149
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1644511149
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_841
timestamp 1644511149
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_853
timestamp 1644511149
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_865
timestamp 1644511149
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_877
timestamp 1644511149
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1644511149
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1644511149
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_897
timestamp 1644511149
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_909
timestamp 1644511149
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_921
timestamp 1644511149
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_933
timestamp 1644511149
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1644511149
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1644511149
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_953
timestamp 1644511149
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_965
timestamp 1644511149
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_977
timestamp 1644511149
transform 1 0 90988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_992
timestamp 1644511149
transform 1 0 92368 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1004
timestamp 1644511149
transform 1 0 93472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1009
timestamp 1644511149
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1021
timestamp 1644511149
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1033
timestamp 1644511149
transform 1 0 96140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1055
timestamp 1644511149
transform 1 0 98164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1644511149
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1065
timestamp 1644511149
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1077
timestamp 1644511149
transform 1 0 100188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1084
timestamp 1644511149
transform 1 0 100832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1096
timestamp 1644511149
transform 1 0 101936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1116
timestamp 1644511149
transform 1 0 103776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1121
timestamp 1644511149
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1133
timestamp 1644511149
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1161
timestamp 1644511149
transform 1 0 107916 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_1173
timestamp 1644511149
transform 1 0 109020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1177
timestamp 1644511149
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1189
timestamp 1644511149
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1201
timestamp 1644511149
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1213
timestamp 1644511149
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1644511149
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1644511149
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1233
timestamp 1644511149
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1245
timestamp 1644511149
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1257
timestamp 1644511149
transform 1 0 116748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1273
timestamp 1644511149
transform 1 0 118220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1644511149
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1644511149
transform 1 0 10120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1644511149
transform 1 0 11224 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_122
timestamp 1644511149
transform 1 0 12328 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1644511149
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_176
timestamp 1644511149
transform 1 0 17296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_713
timestamp 1644511149
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_737
timestamp 1644511149
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1644511149
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1644511149
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_757
timestamp 1644511149
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_769
timestamp 1644511149
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_781
timestamp 1644511149
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_793
timestamp 1644511149
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1644511149
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1644511149
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_829
timestamp 1644511149
transform 1 0 77372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_841
timestamp 1644511149
transform 1 0 78476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_853
timestamp 1644511149
transform 1 0 79580 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_865
timestamp 1644511149
transform 1 0 80684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_869
timestamp 1644511149
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_881
timestamp 1644511149
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_893
timestamp 1644511149
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_905
timestamp 1644511149
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1644511149
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1644511149
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_925
timestamp 1644511149
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_937
timestamp 1644511149
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_949
timestamp 1644511149
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_961
timestamp 1644511149
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1644511149
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1644511149
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_981
timestamp 1644511149
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_993
timestamp 1644511149
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1005
timestamp 1644511149
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1017
timestamp 1644511149
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1644511149
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1644511149
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1037
timestamp 1644511149
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1049
timestamp 1644511149
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1061
timestamp 1644511149
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1073
timestamp 1644511149
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1644511149
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1644511149
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1093
timestamp 1644511149
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1105
timestamp 1644511149
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1117
timestamp 1644511149
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1129
timestamp 1644511149
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1644511149
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1644511149
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1149
timestamp 1644511149
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1161
timestamp 1644511149
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1173
timestamp 1644511149
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1185
timestamp 1644511149
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1644511149
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1644511149
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1205
timestamp 1644511149
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1217
timestamp 1644511149
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1229
timestamp 1644511149
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1241
timestamp 1644511149
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1644511149
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1644511149
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1261
timestamp 1644511149
transform 1 0 117116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_1273
timestamp 1644511149
transform 1 0 118220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1644511149
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1644511149
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1644511149
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_741
timestamp 1644511149
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_753
timestamp 1644511149
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_765
timestamp 1644511149
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1644511149
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1644511149
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_785
timestamp 1644511149
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_797
timestamp 1644511149
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_809
timestamp 1644511149
transform 1 0 75532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_815
timestamp 1644511149
transform 1 0 76084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_830
timestamp 1644511149
transform 1 0 77464 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_838
timestamp 1644511149
transform 1 0 78200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_841
timestamp 1644511149
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_853
timestamp 1644511149
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_865
timestamp 1644511149
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_877
timestamp 1644511149
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1644511149
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1644511149
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_897
timestamp 1644511149
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_909
timestamp 1644511149
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_921
timestamp 1644511149
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_933
timestamp 1644511149
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1644511149
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1644511149
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_953
timestamp 1644511149
transform 1 0 88780 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_965
timestamp 1644511149
transform 1 0 89884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_977
timestamp 1644511149
transform 1 0 90988 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_989
timestamp 1644511149
transform 1 0 92092 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1001
timestamp 1644511149
transform 1 0 93196 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1644511149
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1009
timestamp 1644511149
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1021
timestamp 1644511149
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1033
timestamp 1644511149
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1045
timestamp 1644511149
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1644511149
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1644511149
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1065
timestamp 1644511149
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1077
timestamp 1644511149
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1089
timestamp 1644511149
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1101
timestamp 1644511149
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1644511149
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1644511149
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1121
timestamp 1644511149
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1133
timestamp 1644511149
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1145
timestamp 1644511149
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1157
timestamp 1644511149
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1644511149
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1644511149
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1177
timestamp 1644511149
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1189
timestamp 1644511149
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1201
timestamp 1644511149
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1213
timestamp 1644511149
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1644511149
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1644511149
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1233
timestamp 1644511149
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1245
timestamp 1644511149
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1257
timestamp 1644511149
transform 1 0 116748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1269
timestamp 1644511149
transform 1 0 117852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_725
timestamp 1644511149
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_737
timestamp 1644511149
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1644511149
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1644511149
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_757
timestamp 1644511149
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_769
timestamp 1644511149
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1644511149
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_793
timestamp 1644511149
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1644511149
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1644511149
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_813
timestamp 1644511149
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_825
timestamp 1644511149
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_837
timestamp 1644511149
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_849
timestamp 1644511149
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1644511149
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1644511149
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_869
timestamp 1644511149
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_881
timestamp 1644511149
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_893
timestamp 1644511149
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_905
timestamp 1644511149
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1644511149
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1644511149
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_925
timestamp 1644511149
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_937
timestamp 1644511149
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_949
timestamp 1644511149
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_961
timestamp 1644511149
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1644511149
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1644511149
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_981
timestamp 1644511149
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_993
timestamp 1644511149
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1005
timestamp 1644511149
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1017
timestamp 1644511149
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1644511149
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1644511149
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1037
timestamp 1644511149
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1049
timestamp 1644511149
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1061
timestamp 1644511149
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1073
timestamp 1644511149
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1644511149
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1644511149
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1093
timestamp 1644511149
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1105
timestamp 1644511149
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1117
timestamp 1644511149
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1129
timestamp 1644511149
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1644511149
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1644511149
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1149
timestamp 1644511149
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1161
timestamp 1644511149
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1173
timestamp 1644511149
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1185
timestamp 1644511149
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1644511149
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1644511149
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1205
timestamp 1644511149
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1217
timestamp 1644511149
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1229
timestamp 1644511149
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1241
timestamp 1644511149
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1644511149
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1644511149
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_1261
timestamp 1644511149
transform 1 0 117116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1273
timestamp 1644511149
transform 1 0 118220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_741
timestamp 1644511149
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_753
timestamp 1644511149
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_765
timestamp 1644511149
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1644511149
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1644511149
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_785
timestamp 1644511149
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_797
timestamp 1644511149
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_809
timestamp 1644511149
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_821
timestamp 1644511149
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1644511149
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1644511149
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_841
timestamp 1644511149
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_853
timestamp 1644511149
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_865
timestamp 1644511149
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_877
timestamp 1644511149
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1644511149
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1644511149
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_897
timestamp 1644511149
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_909
timestamp 1644511149
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_921
timestamp 1644511149
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_933
timestamp 1644511149
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1644511149
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1644511149
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_953
timestamp 1644511149
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_965
timestamp 1644511149
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_977
timestamp 1644511149
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_989
timestamp 1644511149
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1644511149
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1644511149
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1009
timestamp 1644511149
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1021
timestamp 1644511149
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1033
timestamp 1644511149
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1045
timestamp 1644511149
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1644511149
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1644511149
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1065
timestamp 1644511149
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1077
timestamp 1644511149
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1089
timestamp 1644511149
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1101
timestamp 1644511149
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1644511149
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1644511149
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1121
timestamp 1644511149
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1133
timestamp 1644511149
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1145
timestamp 1644511149
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1157
timestamp 1644511149
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1644511149
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1644511149
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1177
timestamp 1644511149
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1189
timestamp 1644511149
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1201
timestamp 1644511149
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1213
timestamp 1644511149
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1644511149
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1644511149
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1233
timestamp 1644511149
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1245
timestamp 1644511149
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1257
timestamp 1644511149
transform 1 0 116748 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1269
timestamp 1644511149
transform 1 0 117852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1644511149
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_725
timestamp 1644511149
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_737
timestamp 1644511149
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1644511149
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1644511149
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_757
timestamp 1644511149
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_769
timestamp 1644511149
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_781
timestamp 1644511149
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_793
timestamp 1644511149
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1644511149
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1644511149
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_813
timestamp 1644511149
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_825
timestamp 1644511149
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_837
timestamp 1644511149
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_849
timestamp 1644511149
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1644511149
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1644511149
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_869
timestamp 1644511149
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_881
timestamp 1644511149
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_893
timestamp 1644511149
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_905
timestamp 1644511149
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1644511149
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1644511149
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_925
timestamp 1644511149
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_937
timestamp 1644511149
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_949
timestamp 1644511149
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_961
timestamp 1644511149
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1644511149
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1644511149
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_981
timestamp 1644511149
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_993
timestamp 1644511149
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1005
timestamp 1644511149
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1017
timestamp 1644511149
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1644511149
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1644511149
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1037
timestamp 1644511149
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1049
timestamp 1644511149
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1061
timestamp 1644511149
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1073
timestamp 1644511149
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1644511149
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1644511149
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1093
timestamp 1644511149
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1105
timestamp 1644511149
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1117
timestamp 1644511149
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1129
timestamp 1644511149
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1644511149
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1644511149
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1149
timestamp 1644511149
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1161
timestamp 1644511149
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1173
timestamp 1644511149
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1185
timestamp 1644511149
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1644511149
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1644511149
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1205
timestamp 1644511149
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1217
timestamp 1644511149
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1229
timestamp 1644511149
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1241
timestamp 1644511149
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1644511149
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1644511149
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1261
timestamp 1644511149
transform 1 0 117116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1273
timestamp 1644511149
transform 1 0 118220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_235
timestamp 1644511149
transform 1 0 22724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_247
timestamp 1644511149
transform 1 0 23828 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_259
timestamp 1644511149
transform 1 0 24932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp 1644511149
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_741
timestamp 1644511149
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_753
timestamp 1644511149
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_765
timestamp 1644511149
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1644511149
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1644511149
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_785
timestamp 1644511149
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_797
timestamp 1644511149
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_809
timestamp 1644511149
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_821
timestamp 1644511149
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1644511149
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1644511149
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_841
timestamp 1644511149
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_853
timestamp 1644511149
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_865
timestamp 1644511149
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_877
timestamp 1644511149
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1644511149
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1644511149
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_897
timestamp 1644511149
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_909
timestamp 1644511149
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_921
timestamp 1644511149
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_933
timestamp 1644511149
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1644511149
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1644511149
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_953
timestamp 1644511149
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_965
timestamp 1644511149
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_977
timestamp 1644511149
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_989
timestamp 1644511149
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1644511149
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1644511149
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1009
timestamp 1644511149
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1021
timestamp 1644511149
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1033
timestamp 1644511149
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1045
timestamp 1644511149
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1644511149
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1644511149
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1065
timestamp 1644511149
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1077
timestamp 1644511149
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1089
timestamp 1644511149
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1101
timestamp 1644511149
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1644511149
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1644511149
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1121
timestamp 1644511149
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1133
timestamp 1644511149
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1145
timestamp 1644511149
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1157
timestamp 1644511149
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1644511149
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1644511149
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1177
timestamp 1644511149
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1189
timestamp 1644511149
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1201
timestamp 1644511149
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1213
timestamp 1644511149
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1644511149
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1644511149
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1233
timestamp 1644511149
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1245
timestamp 1644511149
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1257
timestamp 1644511149
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1269
timestamp 1644511149
transform 1 0 117852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_737
timestamp 1644511149
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1644511149
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1644511149
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_757
timestamp 1644511149
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_769
timestamp 1644511149
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_781
timestamp 1644511149
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_793
timestamp 1644511149
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1644511149
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1644511149
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_813
timestamp 1644511149
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_825
timestamp 1644511149
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_837
timestamp 1644511149
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_849
timestamp 1644511149
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1644511149
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1644511149
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_869
timestamp 1644511149
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_881
timestamp 1644511149
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_893
timestamp 1644511149
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_905
timestamp 1644511149
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1644511149
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1644511149
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_925
timestamp 1644511149
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_937
timestamp 1644511149
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_949
timestamp 1644511149
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_961
timestamp 1644511149
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1644511149
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1644511149
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_981
timestamp 1644511149
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_993
timestamp 1644511149
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1005
timestamp 1644511149
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1017
timestamp 1644511149
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1644511149
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1644511149
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1037
timestamp 1644511149
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1049
timestamp 1644511149
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1061
timestamp 1644511149
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1073
timestamp 1644511149
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1644511149
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1644511149
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1093
timestamp 1644511149
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1105
timestamp 1644511149
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1117
timestamp 1644511149
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1129
timestamp 1644511149
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1644511149
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1644511149
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1149
timestamp 1644511149
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1161
timestamp 1644511149
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1173
timestamp 1644511149
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1185
timestamp 1644511149
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1644511149
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1644511149
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1205
timestamp 1644511149
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1217
timestamp 1644511149
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1229
timestamp 1644511149
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1241
timestamp 1644511149
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1644511149
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1644511149
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1261
timestamp 1644511149
transform 1 0 117116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1273
timestamp 1644511149
transform 1 0 118220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_19
timestamp 1644511149
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1644511149
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_741
timestamp 1644511149
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_753
timestamp 1644511149
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_765
timestamp 1644511149
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1644511149
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1644511149
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_785
timestamp 1644511149
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_797
timestamp 1644511149
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_809
timestamp 1644511149
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_821
timestamp 1644511149
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1644511149
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1644511149
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_841
timestamp 1644511149
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_853
timestamp 1644511149
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_865
timestamp 1644511149
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_877
timestamp 1644511149
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1644511149
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1644511149
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_897
timestamp 1644511149
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_909
timestamp 1644511149
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_921
timestamp 1644511149
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_933
timestamp 1644511149
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1644511149
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1644511149
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_953
timestamp 1644511149
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_965
timestamp 1644511149
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_977
timestamp 1644511149
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_989
timestamp 1644511149
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1644511149
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1644511149
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1009
timestamp 1644511149
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1021
timestamp 1644511149
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1033
timestamp 1644511149
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1045
timestamp 1644511149
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1644511149
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1644511149
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1065
timestamp 1644511149
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1077
timestamp 1644511149
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1089
timestamp 1644511149
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1101
timestamp 1644511149
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1644511149
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1644511149
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1121
timestamp 1644511149
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1133
timestamp 1644511149
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1145
timestamp 1644511149
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1157
timestamp 1644511149
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1644511149
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1644511149
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1177
timestamp 1644511149
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1189
timestamp 1644511149
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1201
timestamp 1644511149
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1213
timestamp 1644511149
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1644511149
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1644511149
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1233
timestamp 1644511149
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1245
timestamp 1644511149
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1257
timestamp 1644511149
transform 1 0 116748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1269
timestamp 1644511149
transform 1 0 117852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_737
timestamp 1644511149
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1644511149
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1644511149
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_757
timestamp 1644511149
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_769
timestamp 1644511149
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_781
timestamp 1644511149
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_793
timestamp 1644511149
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1644511149
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1644511149
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_813
timestamp 1644511149
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_825
timestamp 1644511149
transform 1 0 77004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_837
timestamp 1644511149
transform 1 0 78108 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_849
timestamp 1644511149
transform 1 0 79212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_861
timestamp 1644511149
transform 1 0 80316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_867
timestamp 1644511149
transform 1 0 80868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_869
timestamp 1644511149
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_881
timestamp 1644511149
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_893
timestamp 1644511149
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_905
timestamp 1644511149
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1644511149
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1644511149
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_925
timestamp 1644511149
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_937
timestamp 1644511149
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_949
timestamp 1644511149
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_961
timestamp 1644511149
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1644511149
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1644511149
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_981
timestamp 1644511149
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_993
timestamp 1644511149
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1005
timestamp 1644511149
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1017
timestamp 1644511149
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1644511149
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1644511149
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1037
timestamp 1644511149
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1049
timestamp 1644511149
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1061
timestamp 1644511149
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1073
timestamp 1644511149
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1644511149
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1644511149
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1093
timestamp 1644511149
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1105
timestamp 1644511149
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1117
timestamp 1644511149
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1129
timestamp 1644511149
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1644511149
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1644511149
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1149
timestamp 1644511149
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1161
timestamp 1644511149
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1173
timestamp 1644511149
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1185
timestamp 1644511149
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1644511149
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1644511149
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1205
timestamp 1644511149
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1217
timestamp 1644511149
transform 1 0 113068 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1229
timestamp 1644511149
transform 1 0 114172 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1241
timestamp 1644511149
transform 1 0 115276 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1644511149
transform 1 0 116380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1644511149
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1261
timestamp 1644511149
transform 1 0 117116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1273
timestamp 1644511149
transform 1 0 118220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_741
timestamp 1644511149
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_753
timestamp 1644511149
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_765
timestamp 1644511149
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1644511149
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1644511149
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_785
timestamp 1644511149
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_797
timestamp 1644511149
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_809
timestamp 1644511149
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_821
timestamp 1644511149
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1644511149
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1644511149
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_841
timestamp 1644511149
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_853
timestamp 1644511149
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_865
timestamp 1644511149
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_877
timestamp 1644511149
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1644511149
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1644511149
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_897
timestamp 1644511149
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_909
timestamp 1644511149
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_921
timestamp 1644511149
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_933
timestamp 1644511149
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1644511149
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1644511149
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_953
timestamp 1644511149
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_965
timestamp 1644511149
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_977
timestamp 1644511149
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_989
timestamp 1644511149
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1644511149
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1644511149
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1009
timestamp 1644511149
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1021
timestamp 1644511149
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1033
timestamp 1644511149
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1045
timestamp 1644511149
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1644511149
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1644511149
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1065
timestamp 1644511149
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1077
timestamp 1644511149
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1089
timestamp 1644511149
transform 1 0 101292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1101
timestamp 1644511149
transform 1 0 102396 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1113
timestamp 1644511149
transform 1 0 103500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1119
timestamp 1644511149
transform 1 0 104052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1121
timestamp 1644511149
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1133
timestamp 1644511149
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1145
timestamp 1644511149
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1157
timestamp 1644511149
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1644511149
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1644511149
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1177
timestamp 1644511149
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1189
timestamp 1644511149
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1201
timestamp 1644511149
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1213
timestamp 1644511149
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1644511149
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1644511149
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1233
timestamp 1644511149
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1245
timestamp 1644511149
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1257
timestamp 1644511149
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1269
timestamp 1644511149
transform 1 0 117852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1644511149
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_737
timestamp 1644511149
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1644511149
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1644511149
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_757
timestamp 1644511149
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_769
timestamp 1644511149
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_781
timestamp 1644511149
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_793
timestamp 1644511149
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1644511149
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1644511149
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_813
timestamp 1644511149
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_825
timestamp 1644511149
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_837
timestamp 1644511149
transform 1 0 78108 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_849
timestamp 1644511149
transform 1 0 79212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_861
timestamp 1644511149
transform 1 0 80316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_867
timestamp 1644511149
transform 1 0 80868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_869
timestamp 1644511149
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_881
timestamp 1644511149
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_893
timestamp 1644511149
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_905
timestamp 1644511149
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1644511149
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1644511149
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_925
timestamp 1644511149
transform 1 0 86204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_937
timestamp 1644511149
transform 1 0 87308 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_949
timestamp 1644511149
transform 1 0 88412 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_961
timestamp 1644511149
transform 1 0 89516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_973
timestamp 1644511149
transform 1 0 90620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_979
timestamp 1644511149
transform 1 0 91172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_981
timestamp 1644511149
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_993
timestamp 1644511149
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1005
timestamp 1644511149
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1017
timestamp 1644511149
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1644511149
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1644511149
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1037
timestamp 1644511149
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1049
timestamp 1644511149
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1061
timestamp 1644511149
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1073
timestamp 1644511149
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1644511149
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1644511149
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1093
timestamp 1644511149
transform 1 0 101660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1105
timestamp 1644511149
transform 1 0 102764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1117
timestamp 1644511149
transform 1 0 103868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1129
timestamp 1644511149
transform 1 0 104972 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1141
timestamp 1644511149
transform 1 0 106076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1147
timestamp 1644511149
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1149
timestamp 1644511149
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1161
timestamp 1644511149
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1173
timestamp 1644511149
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1185
timestamp 1644511149
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1644511149
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1644511149
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1205
timestamp 1644511149
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1217
timestamp 1644511149
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1229
timestamp 1644511149
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1241
timestamp 1644511149
transform 1 0 115276 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1253
timestamp 1644511149
transform 1 0 116380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1259
timestamp 1644511149
transform 1 0 116932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1261
timestamp 1644511149
transform 1 0 117116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1273
timestamp 1644511149
transform 1 0 118220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_741
timestamp 1644511149
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_753
timestamp 1644511149
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_765
timestamp 1644511149
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1644511149
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1644511149
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_785
timestamp 1644511149
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_797
timestamp 1644511149
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_809
timestamp 1644511149
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_821
timestamp 1644511149
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1644511149
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1644511149
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_841
timestamp 1644511149
transform 1 0 78476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_853
timestamp 1644511149
transform 1 0 79580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_865
timestamp 1644511149
transform 1 0 80684 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_877
timestamp 1644511149
transform 1 0 81788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_889
timestamp 1644511149
transform 1 0 82892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1644511149
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_897
timestamp 1644511149
transform 1 0 83628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_909
timestamp 1644511149
transform 1 0 84732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_921
timestamp 1644511149
transform 1 0 85836 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_933
timestamp 1644511149
transform 1 0 86940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1644511149
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1644511149
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_953
timestamp 1644511149
transform 1 0 88780 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_965
timestamp 1644511149
transform 1 0 89884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_977
timestamp 1644511149
transform 1 0 90988 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_989
timestamp 1644511149
transform 1 0 92092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1644511149
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1644511149
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1009
timestamp 1644511149
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1021
timestamp 1644511149
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1033
timestamp 1644511149
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1045
timestamp 1644511149
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1644511149
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1644511149
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1065
timestamp 1644511149
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1077
timestamp 1644511149
transform 1 0 100188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1089
timestamp 1644511149
transform 1 0 101292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1101
timestamp 1644511149
transform 1 0 102396 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1113
timestamp 1644511149
transform 1 0 103500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1119
timestamp 1644511149
transform 1 0 104052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1121
timestamp 1644511149
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1133
timestamp 1644511149
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1145
timestamp 1644511149
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1157
timestamp 1644511149
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1644511149
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1644511149
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1177
timestamp 1644511149
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1189
timestamp 1644511149
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1201
timestamp 1644511149
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1213
timestamp 1644511149
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1225
timestamp 1644511149
transform 1 0 113804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1231
timestamp 1644511149
transform 1 0 114356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1233
timestamp 1644511149
transform 1 0 114540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1245
timestamp 1644511149
transform 1 0 115644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1257
timestamp 1644511149
transform 1 0 116748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1269
timestamp 1644511149
transform 1 0 117852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_737
timestamp 1644511149
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1644511149
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1644511149
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_757
timestamp 1644511149
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_769
timestamp 1644511149
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_781
timestamp 1644511149
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_793
timestamp 1644511149
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1644511149
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1644511149
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_813
timestamp 1644511149
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_825
timestamp 1644511149
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_837
timestamp 1644511149
transform 1 0 78108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_849
timestamp 1644511149
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1644511149
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1644511149
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_869
timestamp 1644511149
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_881
timestamp 1644511149
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_893
timestamp 1644511149
transform 1 0 83260 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_905
timestamp 1644511149
transform 1 0 84364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_917
timestamp 1644511149
transform 1 0 85468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1644511149
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_925
timestamp 1644511149
transform 1 0 86204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_937
timestamp 1644511149
transform 1 0 87308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_949
timestamp 1644511149
transform 1 0 88412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_961
timestamp 1644511149
transform 1 0 89516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_973
timestamp 1644511149
transform 1 0 90620 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_979
timestamp 1644511149
transform 1 0 91172 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_981
timestamp 1644511149
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_993
timestamp 1644511149
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1005
timestamp 1644511149
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1017
timestamp 1644511149
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1644511149
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1644511149
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1037
timestamp 1644511149
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1049
timestamp 1644511149
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1061
timestamp 1644511149
transform 1 0 98716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1073
timestamp 1644511149
transform 1 0 99820 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1085
timestamp 1644511149
transform 1 0 100924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1091
timestamp 1644511149
transform 1 0 101476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1093
timestamp 1644511149
transform 1 0 101660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1105
timestamp 1644511149
transform 1 0 102764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1117
timestamp 1644511149
transform 1 0 103868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1129
timestamp 1644511149
transform 1 0 104972 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1141
timestamp 1644511149
transform 1 0 106076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1147
timestamp 1644511149
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1149
timestamp 1644511149
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1161
timestamp 1644511149
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1173
timestamp 1644511149
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1185
timestamp 1644511149
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1644511149
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1644511149
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1205
timestamp 1644511149
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1217
timestamp 1644511149
transform 1 0 113068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1229
timestamp 1644511149
transform 1 0 114172 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1241
timestamp 1644511149
transform 1 0 115276 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1253
timestamp 1644511149
transform 1 0 116380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1644511149
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1261
timestamp 1644511149
transform 1 0 117116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1273
timestamp 1644511149
transform 1 0 118220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_741
timestamp 1644511149
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_753
timestamp 1644511149
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_765
timestamp 1644511149
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1644511149
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1644511149
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_785
timestamp 1644511149
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_797
timestamp 1644511149
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_809
timestamp 1644511149
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_821
timestamp 1644511149
transform 1 0 76636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_833
timestamp 1644511149
transform 1 0 77740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1644511149
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_841
timestamp 1644511149
transform 1 0 78476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_853
timestamp 1644511149
transform 1 0 79580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_865
timestamp 1644511149
transform 1 0 80684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_877
timestamp 1644511149
transform 1 0 81788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_889
timestamp 1644511149
transform 1 0 82892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1644511149
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_897
timestamp 1644511149
transform 1 0 83628 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_909
timestamp 1644511149
transform 1 0 84732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_921
timestamp 1644511149
transform 1 0 85836 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_933
timestamp 1644511149
transform 1 0 86940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1644511149
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1644511149
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_953
timestamp 1644511149
transform 1 0 88780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_965
timestamp 1644511149
transform 1 0 89884 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_977
timestamp 1644511149
transform 1 0 90988 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_989
timestamp 1644511149
transform 1 0 92092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1001
timestamp 1644511149
transform 1 0 93196 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1007
timestamp 1644511149
transform 1 0 93748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1009
timestamp 1644511149
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1021
timestamp 1644511149
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1033
timestamp 1644511149
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1045
timestamp 1644511149
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1057
timestamp 1644511149
transform 1 0 98348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1063
timestamp 1644511149
transform 1 0 98900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1065
timestamp 1644511149
transform 1 0 99084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1077
timestamp 1644511149
transform 1 0 100188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1089
timestamp 1644511149
transform 1 0 101292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1101
timestamp 1644511149
transform 1 0 102396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1113
timestamp 1644511149
transform 1 0 103500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1119
timestamp 1644511149
transform 1 0 104052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1121
timestamp 1644511149
transform 1 0 104236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1133
timestamp 1644511149
transform 1 0 105340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1145
timestamp 1644511149
transform 1 0 106444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1157
timestamp 1644511149
transform 1 0 107548 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1169
timestamp 1644511149
transform 1 0 108652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1175
timestamp 1644511149
transform 1 0 109204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1177
timestamp 1644511149
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1189
timestamp 1644511149
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1201
timestamp 1644511149
transform 1 0 111596 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1213
timestamp 1644511149
transform 1 0 112700 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1225
timestamp 1644511149
transform 1 0 113804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1231
timestamp 1644511149
transform 1 0 114356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1233
timestamp 1644511149
transform 1 0 114540 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1245
timestamp 1644511149
transform 1 0 115644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1257
timestamp 1644511149
transform 1 0 116748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1269
timestamp 1644511149
transform 1 0 117852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_725
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_737
timestamp 1644511149
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1644511149
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1644511149
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_757
timestamp 1644511149
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_769
timestamp 1644511149
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_781
timestamp 1644511149
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_793
timestamp 1644511149
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1644511149
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1644511149
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_813
timestamp 1644511149
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_825
timestamp 1644511149
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_837
timestamp 1644511149
transform 1 0 78108 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_849
timestamp 1644511149
transform 1 0 79212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1644511149
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1644511149
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_869
timestamp 1644511149
transform 1 0 81052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_881
timestamp 1644511149
transform 1 0 82156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_893
timestamp 1644511149
transform 1 0 83260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_905
timestamp 1644511149
transform 1 0 84364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_917
timestamp 1644511149
transform 1 0 85468 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1644511149
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_925
timestamp 1644511149
transform 1 0 86204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_937
timestamp 1644511149
transform 1 0 87308 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_949
timestamp 1644511149
transform 1 0 88412 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_961
timestamp 1644511149
transform 1 0 89516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1644511149
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1644511149
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_981
timestamp 1644511149
transform 1 0 91356 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_993
timestamp 1644511149
transform 1 0 92460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1005
timestamp 1644511149
transform 1 0 93564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1017
timestamp 1644511149
transform 1 0 94668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1029
timestamp 1644511149
transform 1 0 95772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1035
timestamp 1644511149
transform 1 0 96324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1037
timestamp 1644511149
transform 1 0 96508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1049
timestamp 1644511149
transform 1 0 97612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1061
timestamp 1644511149
transform 1 0 98716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1073
timestamp 1644511149
transform 1 0 99820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1085
timestamp 1644511149
transform 1 0 100924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1091
timestamp 1644511149
transform 1 0 101476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1093
timestamp 1644511149
transform 1 0 101660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1105
timestamp 1644511149
transform 1 0 102764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1117
timestamp 1644511149
transform 1 0 103868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1129
timestamp 1644511149
transform 1 0 104972 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1644511149
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1644511149
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1149
timestamp 1644511149
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1161
timestamp 1644511149
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1173
timestamp 1644511149
transform 1 0 109020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1185
timestamp 1644511149
transform 1 0 110124 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1197
timestamp 1644511149
transform 1 0 111228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1203
timestamp 1644511149
transform 1 0 111780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1205
timestamp 1644511149
transform 1 0 111964 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1217
timestamp 1644511149
transform 1 0 113068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1229
timestamp 1644511149
transform 1 0 114172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1241
timestamp 1644511149
transform 1 0 115276 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1253
timestamp 1644511149
transform 1 0 116380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1259
timestamp 1644511149
transform 1 0 116932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1261
timestamp 1644511149
transform 1 0 117116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1273
timestamp 1644511149
transform 1 0 118220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_741
timestamp 1644511149
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_753
timestamp 1644511149
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_765
timestamp 1644511149
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1644511149
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1644511149
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_785
timestamp 1644511149
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_797
timestamp 1644511149
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_809
timestamp 1644511149
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_821
timestamp 1644511149
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_833
timestamp 1644511149
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_839
timestamp 1644511149
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_841
timestamp 1644511149
transform 1 0 78476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_853
timestamp 1644511149
transform 1 0 79580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_865
timestamp 1644511149
transform 1 0 80684 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_877
timestamp 1644511149
transform 1 0 81788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_889
timestamp 1644511149
transform 1 0 82892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_895
timestamp 1644511149
transform 1 0 83444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_897
timestamp 1644511149
transform 1 0 83628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_909
timestamp 1644511149
transform 1 0 84732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_921
timestamp 1644511149
transform 1 0 85836 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_933
timestamp 1644511149
transform 1 0 86940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_945
timestamp 1644511149
transform 1 0 88044 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_951
timestamp 1644511149
transform 1 0 88596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_953
timestamp 1644511149
transform 1 0 88780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_965
timestamp 1644511149
transform 1 0 89884 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_977
timestamp 1644511149
transform 1 0 90988 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_989
timestamp 1644511149
transform 1 0 92092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1001
timestamp 1644511149
transform 1 0 93196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1007
timestamp 1644511149
transform 1 0 93748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1009
timestamp 1644511149
transform 1 0 93932 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1021
timestamp 1644511149
transform 1 0 95036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1033
timestamp 1644511149
transform 1 0 96140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1045
timestamp 1644511149
transform 1 0 97244 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1057
timestamp 1644511149
transform 1 0 98348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1063
timestamp 1644511149
transform 1 0 98900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1065
timestamp 1644511149
transform 1 0 99084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1077
timestamp 1644511149
transform 1 0 100188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1089
timestamp 1644511149
transform 1 0 101292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1101
timestamp 1644511149
transform 1 0 102396 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1113
timestamp 1644511149
transform 1 0 103500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1119
timestamp 1644511149
transform 1 0 104052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1121
timestamp 1644511149
transform 1 0 104236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1133
timestamp 1644511149
transform 1 0 105340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1145
timestamp 1644511149
transform 1 0 106444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1157
timestamp 1644511149
transform 1 0 107548 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1169
timestamp 1644511149
transform 1 0 108652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1175
timestamp 1644511149
transform 1 0 109204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1177
timestamp 1644511149
transform 1 0 109388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1189
timestamp 1644511149
transform 1 0 110492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1201
timestamp 1644511149
transform 1 0 111596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1213
timestamp 1644511149
transform 1 0 112700 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1225
timestamp 1644511149
transform 1 0 113804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1231
timestamp 1644511149
transform 1 0 114356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1233
timestamp 1644511149
transform 1 0 114540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1245
timestamp 1644511149
transform 1 0 115644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1257
timestamp 1644511149
transform 1 0 116748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1269
timestamp 1644511149
transform 1 0 117852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1644511149
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_725
timestamp 1644511149
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_737
timestamp 1644511149
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1644511149
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1644511149
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_757
timestamp 1644511149
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_769
timestamp 1644511149
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_781
timestamp 1644511149
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_793
timestamp 1644511149
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1644511149
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1644511149
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_813
timestamp 1644511149
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_825
timestamp 1644511149
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_837
timestamp 1644511149
transform 1 0 78108 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_849
timestamp 1644511149
transform 1 0 79212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1644511149
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1644511149
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_869
timestamp 1644511149
transform 1 0 81052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_881
timestamp 1644511149
transform 1 0 82156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_893
timestamp 1644511149
transform 1 0 83260 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_905
timestamp 1644511149
transform 1 0 84364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_917
timestamp 1644511149
transform 1 0 85468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_923
timestamp 1644511149
transform 1 0 86020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_925
timestamp 1644511149
transform 1 0 86204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_937
timestamp 1644511149
transform 1 0 87308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_949
timestamp 1644511149
transform 1 0 88412 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_961
timestamp 1644511149
transform 1 0 89516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_973
timestamp 1644511149
transform 1 0 90620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_979
timestamp 1644511149
transform 1 0 91172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_981
timestamp 1644511149
transform 1 0 91356 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_993
timestamp 1644511149
transform 1 0 92460 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1005
timestamp 1644511149
transform 1 0 93564 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1017
timestamp 1644511149
transform 1 0 94668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1029
timestamp 1644511149
transform 1 0 95772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1035
timestamp 1644511149
transform 1 0 96324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1037
timestamp 1644511149
transform 1 0 96508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1049
timestamp 1644511149
transform 1 0 97612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1061
timestamp 1644511149
transform 1 0 98716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1073
timestamp 1644511149
transform 1 0 99820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1085
timestamp 1644511149
transform 1 0 100924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1091
timestamp 1644511149
transform 1 0 101476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1093
timestamp 1644511149
transform 1 0 101660 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1105
timestamp 1644511149
transform 1 0 102764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1117
timestamp 1644511149
transform 1 0 103868 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1129
timestamp 1644511149
transform 1 0 104972 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1141
timestamp 1644511149
transform 1 0 106076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1147
timestamp 1644511149
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1149
timestamp 1644511149
transform 1 0 106812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1161
timestamp 1644511149
transform 1 0 107916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1173
timestamp 1644511149
transform 1 0 109020 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1185
timestamp 1644511149
transform 1 0 110124 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1197
timestamp 1644511149
transform 1 0 111228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1203
timestamp 1644511149
transform 1 0 111780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1205
timestamp 1644511149
transform 1 0 111964 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1217
timestamp 1644511149
transform 1 0 113068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1229
timestamp 1644511149
transform 1 0 114172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1241
timestamp 1644511149
transform 1 0 115276 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1253
timestamp 1644511149
transform 1 0 116380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1259
timestamp 1644511149
transform 1 0 116932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1261
timestamp 1644511149
transform 1 0 117116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_1273
timestamp 1644511149
transform 1 0 118220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_673
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1644511149
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_697
timestamp 1644511149
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_709
timestamp 1644511149
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1644511149
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1644511149
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_741
timestamp 1644511149
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_753
timestamp 1644511149
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_765
timestamp 1644511149
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1644511149
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1644511149
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_785
timestamp 1644511149
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_797
timestamp 1644511149
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_809
timestamp 1644511149
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_821
timestamp 1644511149
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1644511149
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1644511149
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_841
timestamp 1644511149
transform 1 0 78476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_853
timestamp 1644511149
transform 1 0 79580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_865
timestamp 1644511149
transform 1 0 80684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_877
timestamp 1644511149
transform 1 0 81788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_889
timestamp 1644511149
transform 1 0 82892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_895
timestamp 1644511149
transform 1 0 83444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_897
timestamp 1644511149
transform 1 0 83628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_909
timestamp 1644511149
transform 1 0 84732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_921
timestamp 1644511149
transform 1 0 85836 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_933
timestamp 1644511149
transform 1 0 86940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_945
timestamp 1644511149
transform 1 0 88044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_951
timestamp 1644511149
transform 1 0 88596 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_953
timestamp 1644511149
transform 1 0 88780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_965
timestamp 1644511149
transform 1 0 89884 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_977
timestamp 1644511149
transform 1 0 90988 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_989
timestamp 1644511149
transform 1 0 92092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1001
timestamp 1644511149
transform 1 0 93196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1007
timestamp 1644511149
transform 1 0 93748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1009
timestamp 1644511149
transform 1 0 93932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1021
timestamp 1644511149
transform 1 0 95036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1033
timestamp 1644511149
transform 1 0 96140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1045
timestamp 1644511149
transform 1 0 97244 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1057
timestamp 1644511149
transform 1 0 98348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1063
timestamp 1644511149
transform 1 0 98900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1065
timestamp 1644511149
transform 1 0 99084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1077
timestamp 1644511149
transform 1 0 100188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1089
timestamp 1644511149
transform 1 0 101292 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1101
timestamp 1644511149
transform 1 0 102396 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1113
timestamp 1644511149
transform 1 0 103500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1119
timestamp 1644511149
transform 1 0 104052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1121
timestamp 1644511149
transform 1 0 104236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1133
timestamp 1644511149
transform 1 0 105340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1145
timestamp 1644511149
transform 1 0 106444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1157
timestamp 1644511149
transform 1 0 107548 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1169
timestamp 1644511149
transform 1 0 108652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1175
timestamp 1644511149
transform 1 0 109204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1177
timestamp 1644511149
transform 1 0 109388 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1189
timestamp 1644511149
transform 1 0 110492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1201
timestamp 1644511149
transform 1 0 111596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1213
timestamp 1644511149
transform 1 0 112700 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1225
timestamp 1644511149
transform 1 0 113804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1231
timestamp 1644511149
transform 1 0 114356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1233
timestamp 1644511149
transform 1 0 114540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1245
timestamp 1644511149
transform 1 0 115644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1257
timestamp 1644511149
transform 1 0 116748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1269
timestamp 1644511149
transform 1 0 117852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1644511149
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1644511149
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1644511149
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_737
timestamp 1644511149
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1644511149
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1644511149
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_757
timestamp 1644511149
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_769
timestamp 1644511149
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_781
timestamp 1644511149
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_793
timestamp 1644511149
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1644511149
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1644511149
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_813
timestamp 1644511149
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_825
timestamp 1644511149
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_837
timestamp 1644511149
transform 1 0 78108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_849
timestamp 1644511149
transform 1 0 79212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1644511149
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1644511149
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_869
timestamp 1644511149
transform 1 0 81052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_881
timestamp 1644511149
transform 1 0 82156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_893
timestamp 1644511149
transform 1 0 83260 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_905
timestamp 1644511149
transform 1 0 84364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_917
timestamp 1644511149
transform 1 0 85468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1644511149
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_925
timestamp 1644511149
transform 1 0 86204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_937
timestamp 1644511149
transform 1 0 87308 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_949
timestamp 1644511149
transform 1 0 88412 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_961
timestamp 1644511149
transform 1 0 89516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_973
timestamp 1644511149
transform 1 0 90620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_979
timestamp 1644511149
transform 1 0 91172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_981
timestamp 1644511149
transform 1 0 91356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_993
timestamp 1644511149
transform 1 0 92460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1005
timestamp 1644511149
transform 1 0 93564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1017
timestamp 1644511149
transform 1 0 94668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1029
timestamp 1644511149
transform 1 0 95772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1035
timestamp 1644511149
transform 1 0 96324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1037
timestamp 1644511149
transform 1 0 96508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1049
timestamp 1644511149
transform 1 0 97612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1061
timestamp 1644511149
transform 1 0 98716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1073
timestamp 1644511149
transform 1 0 99820 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1085
timestamp 1644511149
transform 1 0 100924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1091
timestamp 1644511149
transform 1 0 101476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1093
timestamp 1644511149
transform 1 0 101660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1105
timestamp 1644511149
transform 1 0 102764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1117
timestamp 1644511149
transform 1 0 103868 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1129
timestamp 1644511149
transform 1 0 104972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1141
timestamp 1644511149
transform 1 0 106076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1147
timestamp 1644511149
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1149
timestamp 1644511149
transform 1 0 106812 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1161
timestamp 1644511149
transform 1 0 107916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1173
timestamp 1644511149
transform 1 0 109020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1185
timestamp 1644511149
transform 1 0 110124 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1197
timestamp 1644511149
transform 1 0 111228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1203
timestamp 1644511149
transform 1 0 111780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1205
timestamp 1644511149
transform 1 0 111964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1217
timestamp 1644511149
transform 1 0 113068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1229
timestamp 1644511149
transform 1 0 114172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1241
timestamp 1644511149
transform 1 0 115276 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1253
timestamp 1644511149
transform 1 0 116380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1259
timestamp 1644511149
transform 1 0 116932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1261
timestamp 1644511149
transform 1 0 117116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_1273
timestamp 1644511149
transform 1 0 118220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_741
timestamp 1644511149
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_753
timestamp 1644511149
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_765
timestamp 1644511149
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1644511149
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1644511149
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_785
timestamp 1644511149
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_797
timestamp 1644511149
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_809
timestamp 1644511149
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_821
timestamp 1644511149
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1644511149
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1644511149
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_841
timestamp 1644511149
transform 1 0 78476 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_853
timestamp 1644511149
transform 1 0 79580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_865
timestamp 1644511149
transform 1 0 80684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_877
timestamp 1644511149
transform 1 0 81788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_889
timestamp 1644511149
transform 1 0 82892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_895
timestamp 1644511149
transform 1 0 83444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_897
timestamp 1644511149
transform 1 0 83628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_909
timestamp 1644511149
transform 1 0 84732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_921
timestamp 1644511149
transform 1 0 85836 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_933
timestamp 1644511149
transform 1 0 86940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_945
timestamp 1644511149
transform 1 0 88044 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_951
timestamp 1644511149
transform 1 0 88596 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_953
timestamp 1644511149
transform 1 0 88780 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_965
timestamp 1644511149
transform 1 0 89884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_977
timestamp 1644511149
transform 1 0 90988 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_989
timestamp 1644511149
transform 1 0 92092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1001
timestamp 1644511149
transform 1 0 93196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1007
timestamp 1644511149
transform 1 0 93748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1009
timestamp 1644511149
transform 1 0 93932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1021
timestamp 1644511149
transform 1 0 95036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1033
timestamp 1644511149
transform 1 0 96140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1045
timestamp 1644511149
transform 1 0 97244 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1057
timestamp 1644511149
transform 1 0 98348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1063
timestamp 1644511149
transform 1 0 98900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1065
timestamp 1644511149
transform 1 0 99084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1077
timestamp 1644511149
transform 1 0 100188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1089
timestamp 1644511149
transform 1 0 101292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1101
timestamp 1644511149
transform 1 0 102396 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1113
timestamp 1644511149
transform 1 0 103500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1119
timestamp 1644511149
transform 1 0 104052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1121
timestamp 1644511149
transform 1 0 104236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1133
timestamp 1644511149
transform 1 0 105340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1145
timestamp 1644511149
transform 1 0 106444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1157
timestamp 1644511149
transform 1 0 107548 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1169
timestamp 1644511149
transform 1 0 108652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1175
timestamp 1644511149
transform 1 0 109204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1177
timestamp 1644511149
transform 1 0 109388 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1189
timestamp 1644511149
transform 1 0 110492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1201
timestamp 1644511149
transform 1 0 111596 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1213
timestamp 1644511149
transform 1 0 112700 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1225
timestamp 1644511149
transform 1 0 113804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1231
timestamp 1644511149
transform 1 0 114356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1233
timestamp 1644511149
transform 1 0 114540 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1245
timestamp 1644511149
transform 1 0 115644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1257
timestamp 1644511149
transform 1 0 116748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1269
timestamp 1644511149
transform 1 0 117852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_737
timestamp 1644511149
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1644511149
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1644511149
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_757
timestamp 1644511149
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_769
timestamp 1644511149
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_781
timestamp 1644511149
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_793
timestamp 1644511149
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1644511149
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1644511149
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_813
timestamp 1644511149
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_825
timestamp 1644511149
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_837
timestamp 1644511149
transform 1 0 78108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_849
timestamp 1644511149
transform 1 0 79212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_861
timestamp 1644511149
transform 1 0 80316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_867
timestamp 1644511149
transform 1 0 80868 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_869
timestamp 1644511149
transform 1 0 81052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_881
timestamp 1644511149
transform 1 0 82156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_893
timestamp 1644511149
transform 1 0 83260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_905
timestamp 1644511149
transform 1 0 84364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_917
timestamp 1644511149
transform 1 0 85468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_923
timestamp 1644511149
transform 1 0 86020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_925
timestamp 1644511149
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_937
timestamp 1644511149
transform 1 0 87308 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_949
timestamp 1644511149
transform 1 0 88412 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_961
timestamp 1644511149
transform 1 0 89516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_973
timestamp 1644511149
transform 1 0 90620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_979
timestamp 1644511149
transform 1 0 91172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_981
timestamp 1644511149
transform 1 0 91356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_993
timestamp 1644511149
transform 1 0 92460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1005
timestamp 1644511149
transform 1 0 93564 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1017
timestamp 1644511149
transform 1 0 94668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1029
timestamp 1644511149
transform 1 0 95772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1035
timestamp 1644511149
transform 1 0 96324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1037
timestamp 1644511149
transform 1 0 96508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1049
timestamp 1644511149
transform 1 0 97612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1061
timestamp 1644511149
transform 1 0 98716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1073
timestamp 1644511149
transform 1 0 99820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1085
timestamp 1644511149
transform 1 0 100924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1091
timestamp 1644511149
transform 1 0 101476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1093
timestamp 1644511149
transform 1 0 101660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1105
timestamp 1644511149
transform 1 0 102764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1117
timestamp 1644511149
transform 1 0 103868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1129
timestamp 1644511149
transform 1 0 104972 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1141
timestamp 1644511149
transform 1 0 106076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1147
timestamp 1644511149
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1149
timestamp 1644511149
transform 1 0 106812 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1161
timestamp 1644511149
transform 1 0 107916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1173
timestamp 1644511149
transform 1 0 109020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1185
timestamp 1644511149
transform 1 0 110124 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1197
timestamp 1644511149
transform 1 0 111228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1203
timestamp 1644511149
transform 1 0 111780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1205
timestamp 1644511149
transform 1 0 111964 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1217
timestamp 1644511149
transform 1 0 113068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1229
timestamp 1644511149
transform 1 0 114172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1241
timestamp 1644511149
transform 1 0 115276 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1253
timestamp 1644511149
transform 1 0 116380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1259
timestamp 1644511149
transform 1 0 116932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1261
timestamp 1644511149
transform 1 0 117116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_1273
timestamp 1644511149
transform 1 0 118220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_641
timestamp 1644511149
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_653
timestamp 1644511149
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1644511149
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1644511149
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1644511149
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1644511149
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1644511149
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_741
timestamp 1644511149
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_753
timestamp 1644511149
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_765
timestamp 1644511149
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1644511149
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1644511149
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_785
timestamp 1644511149
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_797
timestamp 1644511149
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_809
timestamp 1644511149
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_821
timestamp 1644511149
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1644511149
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1644511149
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_841
timestamp 1644511149
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_853
timestamp 1644511149
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_865
timestamp 1644511149
transform 1 0 80684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_877
timestamp 1644511149
transform 1 0 81788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_889
timestamp 1644511149
transform 1 0 82892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_895
timestamp 1644511149
transform 1 0 83444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_897
timestamp 1644511149
transform 1 0 83628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_909
timestamp 1644511149
transform 1 0 84732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_921
timestamp 1644511149
transform 1 0 85836 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_933
timestamp 1644511149
transform 1 0 86940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_945
timestamp 1644511149
transform 1 0 88044 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_951
timestamp 1644511149
transform 1 0 88596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_953
timestamp 1644511149
transform 1 0 88780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_965
timestamp 1644511149
transform 1 0 89884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_977
timestamp 1644511149
transform 1 0 90988 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_989
timestamp 1644511149
transform 1 0 92092 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1001
timestamp 1644511149
transform 1 0 93196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1007
timestamp 1644511149
transform 1 0 93748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1009
timestamp 1644511149
transform 1 0 93932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1021
timestamp 1644511149
transform 1 0 95036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1033
timestamp 1644511149
transform 1 0 96140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1045
timestamp 1644511149
transform 1 0 97244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1057
timestamp 1644511149
transform 1 0 98348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1063
timestamp 1644511149
transform 1 0 98900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1065
timestamp 1644511149
transform 1 0 99084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1077
timestamp 1644511149
transform 1 0 100188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1089
timestamp 1644511149
transform 1 0 101292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1101
timestamp 1644511149
transform 1 0 102396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1113
timestamp 1644511149
transform 1 0 103500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1119
timestamp 1644511149
transform 1 0 104052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1121
timestamp 1644511149
transform 1 0 104236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1133
timestamp 1644511149
transform 1 0 105340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1145
timestamp 1644511149
transform 1 0 106444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1157
timestamp 1644511149
transform 1 0 107548 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1169
timestamp 1644511149
transform 1 0 108652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1175
timestamp 1644511149
transform 1 0 109204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1177
timestamp 1644511149
transform 1 0 109388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1189
timestamp 1644511149
transform 1 0 110492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1201
timestamp 1644511149
transform 1 0 111596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1213
timestamp 1644511149
transform 1 0 112700 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1225
timestamp 1644511149
transform 1 0 113804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1231
timestamp 1644511149
transform 1 0 114356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1233
timestamp 1644511149
transform 1 0 114540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1245
timestamp 1644511149
transform 1 0 115644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1257
timestamp 1644511149
transform 1 0 116748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1269
timestamp 1644511149
transform 1 0 117852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1644511149
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_725
timestamp 1644511149
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_737
timestamp 1644511149
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1644511149
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1644511149
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_757
timestamp 1644511149
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_769
timestamp 1644511149
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_781
timestamp 1644511149
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_793
timestamp 1644511149
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1644511149
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1644511149
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_813
timestamp 1644511149
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_825
timestamp 1644511149
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_837
timestamp 1644511149
transform 1 0 78108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_849
timestamp 1644511149
transform 1 0 79212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_861
timestamp 1644511149
transform 1 0 80316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_867
timestamp 1644511149
transform 1 0 80868 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_869
timestamp 1644511149
transform 1 0 81052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_881
timestamp 1644511149
transform 1 0 82156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_893
timestamp 1644511149
transform 1 0 83260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_905
timestamp 1644511149
transform 1 0 84364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_917
timestamp 1644511149
transform 1 0 85468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_923
timestamp 1644511149
transform 1 0 86020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_925
timestamp 1644511149
transform 1 0 86204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_937
timestamp 1644511149
transform 1 0 87308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_949
timestamp 1644511149
transform 1 0 88412 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_961
timestamp 1644511149
transform 1 0 89516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_973
timestamp 1644511149
transform 1 0 90620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_979
timestamp 1644511149
transform 1 0 91172 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_981
timestamp 1644511149
transform 1 0 91356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_993
timestamp 1644511149
transform 1 0 92460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1005
timestamp 1644511149
transform 1 0 93564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1017
timestamp 1644511149
transform 1 0 94668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1029
timestamp 1644511149
transform 1 0 95772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1035
timestamp 1644511149
transform 1 0 96324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1037
timestamp 1644511149
transform 1 0 96508 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1049
timestamp 1644511149
transform 1 0 97612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1061
timestamp 1644511149
transform 1 0 98716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1073
timestamp 1644511149
transform 1 0 99820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1085
timestamp 1644511149
transform 1 0 100924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1091
timestamp 1644511149
transform 1 0 101476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1093
timestamp 1644511149
transform 1 0 101660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1105
timestamp 1644511149
transform 1 0 102764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1117
timestamp 1644511149
transform 1 0 103868 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1129
timestamp 1644511149
transform 1 0 104972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1141
timestamp 1644511149
transform 1 0 106076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1147
timestamp 1644511149
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1149
timestamp 1644511149
transform 1 0 106812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1161
timestamp 1644511149
transform 1 0 107916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1173
timestamp 1644511149
transform 1 0 109020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1185
timestamp 1644511149
transform 1 0 110124 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1197
timestamp 1644511149
transform 1 0 111228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1203
timestamp 1644511149
transform 1 0 111780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1205
timestamp 1644511149
transform 1 0 111964 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1217
timestamp 1644511149
transform 1 0 113068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1229
timestamp 1644511149
transform 1 0 114172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1241
timestamp 1644511149
transform 1 0 115276 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1253
timestamp 1644511149
transform 1 0 116380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1259
timestamp 1644511149
transform 1 0 116932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1261
timestamp 1644511149
transform 1 0 117116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_1273
timestamp 1644511149
transform 1 0 118220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_741
timestamp 1644511149
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_753
timestamp 1644511149
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_765
timestamp 1644511149
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1644511149
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1644511149
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_785
timestamp 1644511149
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_797
timestamp 1644511149
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_809
timestamp 1644511149
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_821
timestamp 1644511149
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1644511149
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1644511149
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_841
timestamp 1644511149
transform 1 0 78476 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_853
timestamp 1644511149
transform 1 0 79580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_865
timestamp 1644511149
transform 1 0 80684 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_877
timestamp 1644511149
transform 1 0 81788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_889
timestamp 1644511149
transform 1 0 82892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_895
timestamp 1644511149
transform 1 0 83444 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_897
timestamp 1644511149
transform 1 0 83628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_909
timestamp 1644511149
transform 1 0 84732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_921
timestamp 1644511149
transform 1 0 85836 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_933
timestamp 1644511149
transform 1 0 86940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_945
timestamp 1644511149
transform 1 0 88044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_951
timestamp 1644511149
transform 1 0 88596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_953
timestamp 1644511149
transform 1 0 88780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_965
timestamp 1644511149
transform 1 0 89884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_977
timestamp 1644511149
transform 1 0 90988 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_989
timestamp 1644511149
transform 1 0 92092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1001
timestamp 1644511149
transform 1 0 93196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1007
timestamp 1644511149
transform 1 0 93748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1009
timestamp 1644511149
transform 1 0 93932 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1021
timestamp 1644511149
transform 1 0 95036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1033
timestamp 1644511149
transform 1 0 96140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1045
timestamp 1644511149
transform 1 0 97244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1057
timestamp 1644511149
transform 1 0 98348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1063
timestamp 1644511149
transform 1 0 98900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1065
timestamp 1644511149
transform 1 0 99084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1077
timestamp 1644511149
transform 1 0 100188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1089
timestamp 1644511149
transform 1 0 101292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1101
timestamp 1644511149
transform 1 0 102396 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1113
timestamp 1644511149
transform 1 0 103500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1119
timestamp 1644511149
transform 1 0 104052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1121
timestamp 1644511149
transform 1 0 104236 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1133
timestamp 1644511149
transform 1 0 105340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1145
timestamp 1644511149
transform 1 0 106444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1157
timestamp 1644511149
transform 1 0 107548 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1169
timestamp 1644511149
transform 1 0 108652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1175
timestamp 1644511149
transform 1 0 109204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1177
timestamp 1644511149
transform 1 0 109388 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1189
timestamp 1644511149
transform 1 0 110492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1201
timestamp 1644511149
transform 1 0 111596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1213
timestamp 1644511149
transform 1 0 112700 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1225
timestamp 1644511149
transform 1 0 113804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1231
timestamp 1644511149
transform 1 0 114356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1233
timestamp 1644511149
transform 1 0 114540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1245
timestamp 1644511149
transform 1 0 115644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1257
timestamp 1644511149
transform 1 0 116748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1265
timestamp 1644511149
transform 1 0 117484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_1273
timestamp 1644511149
transform 1 0 118220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_609
timestamp 1644511149
transform 1 0 57132 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_616
timestamp 1644511149
transform 1 0 57776 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_628
timestamp 1644511149
transform 1 0 58880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_640
timestamp 1644511149
transform 1 0 59984 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_725
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_737
timestamp 1644511149
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1644511149
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1644511149
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_757
timestamp 1644511149
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_769
timestamp 1644511149
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_781
timestamp 1644511149
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_793
timestamp 1644511149
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1644511149
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1644511149
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_813
timestamp 1644511149
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_825
timestamp 1644511149
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_837
timestamp 1644511149
transform 1 0 78108 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_849
timestamp 1644511149
transform 1 0 79212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_861
timestamp 1644511149
transform 1 0 80316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_867
timestamp 1644511149
transform 1 0 80868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_869
timestamp 1644511149
transform 1 0 81052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_881
timestamp 1644511149
transform 1 0 82156 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_893
timestamp 1644511149
transform 1 0 83260 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_905
timestamp 1644511149
transform 1 0 84364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_917
timestamp 1644511149
transform 1 0 85468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_923
timestamp 1644511149
transform 1 0 86020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_925
timestamp 1644511149
transform 1 0 86204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_937
timestamp 1644511149
transform 1 0 87308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_949
timestamp 1644511149
transform 1 0 88412 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_961
timestamp 1644511149
transform 1 0 89516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_973
timestamp 1644511149
transform 1 0 90620 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_979
timestamp 1644511149
transform 1 0 91172 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_981
timestamp 1644511149
transform 1 0 91356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_993
timestamp 1644511149
transform 1 0 92460 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1005
timestamp 1644511149
transform 1 0 93564 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1017
timestamp 1644511149
transform 1 0 94668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1029
timestamp 1644511149
transform 1 0 95772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1035
timestamp 1644511149
transform 1 0 96324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1037
timestamp 1644511149
transform 1 0 96508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1049
timestamp 1644511149
transform 1 0 97612 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1061
timestamp 1644511149
transform 1 0 98716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1073
timestamp 1644511149
transform 1 0 99820 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1085
timestamp 1644511149
transform 1 0 100924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1091
timestamp 1644511149
transform 1 0 101476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1093
timestamp 1644511149
transform 1 0 101660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1105
timestamp 1644511149
transform 1 0 102764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1117
timestamp 1644511149
transform 1 0 103868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1129
timestamp 1644511149
transform 1 0 104972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1141
timestamp 1644511149
transform 1 0 106076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1147
timestamp 1644511149
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1149
timestamp 1644511149
transform 1 0 106812 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1161
timestamp 1644511149
transform 1 0 107916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1173
timestamp 1644511149
transform 1 0 109020 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1185
timestamp 1644511149
transform 1 0 110124 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1197
timestamp 1644511149
transform 1 0 111228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1203
timestamp 1644511149
transform 1 0 111780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1205
timestamp 1644511149
transform 1 0 111964 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1217
timestamp 1644511149
transform 1 0 113068 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1229
timestamp 1644511149
transform 1 0 114172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1241
timestamp 1644511149
transform 1 0 115276 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1253
timestamp 1644511149
transform 1 0 116380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1259
timestamp 1644511149
transform 1 0 116932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1261
timestamp 1644511149
transform 1 0 117116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_1273
timestamp 1644511149
transform 1 0 118220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_9
timestamp 1644511149
transform 1 0 1932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_21
timestamp 1644511149
transform 1 0 3036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_33
timestamp 1644511149
transform 1 0 4140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_45
timestamp 1644511149
transform 1 0 5244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_689
timestamp 1644511149
transform 1 0 64492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_710
timestamp 1644511149
transform 1 0 66424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_717
timestamp 1644511149
transform 1 0 67068 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_725
timestamp 1644511149
transform 1 0 67804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_747
timestamp 1644511149
transform 1 0 69828 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_755
timestamp 1644511149
transform 1 0 70564 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_763
timestamp 1644511149
transform 1 0 71300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_775
timestamp 1644511149
transform 1 0 72404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1644511149
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_785
timestamp 1644511149
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_797
timestamp 1644511149
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_809
timestamp 1644511149
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_821
timestamp 1644511149
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1644511149
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1644511149
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_841
timestamp 1644511149
transform 1 0 78476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_853
timestamp 1644511149
transform 1 0 79580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_865
timestamp 1644511149
transform 1 0 80684 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_877
timestamp 1644511149
transform 1 0 81788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_889
timestamp 1644511149
transform 1 0 82892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_895
timestamp 1644511149
transform 1 0 83444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_897
timestamp 1644511149
transform 1 0 83628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_909
timestamp 1644511149
transform 1 0 84732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_921
timestamp 1644511149
transform 1 0 85836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_933
timestamp 1644511149
transform 1 0 86940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_945
timestamp 1644511149
transform 1 0 88044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_951
timestamp 1644511149
transform 1 0 88596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_953
timestamp 1644511149
transform 1 0 88780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_965
timestamp 1644511149
transform 1 0 89884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_977
timestamp 1644511149
transform 1 0 90988 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_989
timestamp 1644511149
transform 1 0 92092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1001
timestamp 1644511149
transform 1 0 93196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1007
timestamp 1644511149
transform 1 0 93748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1009
timestamp 1644511149
transform 1 0 93932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1021
timestamp 1644511149
transform 1 0 95036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1033
timestamp 1644511149
transform 1 0 96140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1045
timestamp 1644511149
transform 1 0 97244 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1057
timestamp 1644511149
transform 1 0 98348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1063
timestamp 1644511149
transform 1 0 98900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1065
timestamp 1644511149
transform 1 0 99084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1077
timestamp 1644511149
transform 1 0 100188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1089
timestamp 1644511149
transform 1 0 101292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1101
timestamp 1644511149
transform 1 0 102396 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1113
timestamp 1644511149
transform 1 0 103500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1119
timestamp 1644511149
transform 1 0 104052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1121
timestamp 1644511149
transform 1 0 104236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1133
timestamp 1644511149
transform 1 0 105340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1145
timestamp 1644511149
transform 1 0 106444 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1157
timestamp 1644511149
transform 1 0 107548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1169
timestamp 1644511149
transform 1 0 108652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1175
timestamp 1644511149
transform 1 0 109204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1177
timestamp 1644511149
transform 1 0 109388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1189
timestamp 1644511149
transform 1 0 110492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1201
timestamp 1644511149
transform 1 0 111596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1213
timestamp 1644511149
transform 1 0 112700 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1225
timestamp 1644511149
transform 1 0 113804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1231
timestamp 1644511149
transform 1 0 114356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1233
timestamp 1644511149
transform 1 0 114540 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1245
timestamp 1644511149
transform 1 0 115644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1257
timestamp 1644511149
transform 1 0 116748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_1273
timestamp 1644511149
transform 1 0 118220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_677
timestamp 1644511149
transform 1 0 63388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_695
timestamp 1644511149
transform 1 0 65044 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_733
timestamp 1644511149
transform 1 0 68540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_739
timestamp 1644511149
transform 1 0 69092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_751
timestamp 1644511149
transform 1 0 70196 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1644511149
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_757
timestamp 1644511149
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_769
timestamp 1644511149
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_781
timestamp 1644511149
transform 1 0 72956 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_803
timestamp 1644511149
transform 1 0 74980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1644511149
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_813
timestamp 1644511149
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_825
timestamp 1644511149
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_837
timestamp 1644511149
transform 1 0 78108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_849
timestamp 1644511149
transform 1 0 79212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_861
timestamp 1644511149
transform 1 0 80316 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_867
timestamp 1644511149
transform 1 0 80868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_869
timestamp 1644511149
transform 1 0 81052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_881
timestamp 1644511149
transform 1 0 82156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_893
timestamp 1644511149
transform 1 0 83260 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_905
timestamp 1644511149
transform 1 0 84364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_917
timestamp 1644511149
transform 1 0 85468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_923
timestamp 1644511149
transform 1 0 86020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_925
timestamp 1644511149
transform 1 0 86204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_937
timestamp 1644511149
transform 1 0 87308 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_949
timestamp 1644511149
transform 1 0 88412 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_961
timestamp 1644511149
transform 1 0 89516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_973
timestamp 1644511149
transform 1 0 90620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_979
timestamp 1644511149
transform 1 0 91172 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_981
timestamp 1644511149
transform 1 0 91356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_993
timestamp 1644511149
transform 1 0 92460 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1005
timestamp 1644511149
transform 1 0 93564 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1017
timestamp 1644511149
transform 1 0 94668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1029
timestamp 1644511149
transform 1 0 95772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1035
timestamp 1644511149
transform 1 0 96324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1037
timestamp 1644511149
transform 1 0 96508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1049
timestamp 1644511149
transform 1 0 97612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1061
timestamp 1644511149
transform 1 0 98716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1073
timestamp 1644511149
transform 1 0 99820 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1085
timestamp 1644511149
transform 1 0 100924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1091
timestamp 1644511149
transform 1 0 101476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1093
timestamp 1644511149
transform 1 0 101660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1105
timestamp 1644511149
transform 1 0 102764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1117
timestamp 1644511149
transform 1 0 103868 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1129
timestamp 1644511149
transform 1 0 104972 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1141
timestamp 1644511149
transform 1 0 106076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1147
timestamp 1644511149
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1149
timestamp 1644511149
transform 1 0 106812 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1161
timestamp 1644511149
transform 1 0 107916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1173
timestamp 1644511149
transform 1 0 109020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1185
timestamp 1644511149
transform 1 0 110124 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1197
timestamp 1644511149
transform 1 0 111228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1203
timestamp 1644511149
transform 1 0 111780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1205
timestamp 1644511149
transform 1 0 111964 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1217
timestamp 1644511149
transform 1 0 113068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1229
timestamp 1644511149
transform 1 0 114172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1241
timestamp 1644511149
transform 1 0 115276 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1253
timestamp 1644511149
transform 1 0 116380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1259
timestamp 1644511149
transform 1 0 116932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1261
timestamp 1644511149
transform 1 0 117116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1273
timestamp 1644511149
transform 1 0 118220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1644511149
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_673
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_685
timestamp 1644511149
transform 1 0 64124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_693
timestamp 1644511149
transform 1 0 64860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_697
timestamp 1644511149
transform 1 0 65228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_708
timestamp 1644511149
transform 1 0 66240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_720
timestamp 1644511149
transform 1 0 67344 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_738
timestamp 1644511149
transform 1 0 69000 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_758
timestamp 1644511149
transform 1 0 70840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_770
timestamp 1644511149
transform 1 0 71944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_782
timestamp 1644511149
transform 1 0 73048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_785
timestamp 1644511149
transform 1 0 73324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_790
timestamp 1644511149
transform 1 0 73784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_803
timestamp 1644511149
transform 1 0 74980 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_815
timestamp 1644511149
transform 1 0 76084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_827
timestamp 1644511149
transform 1 0 77188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1644511149
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_841
timestamp 1644511149
transform 1 0 78476 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_853
timestamp 1644511149
transform 1 0 79580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_865
timestamp 1644511149
transform 1 0 80684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_877
timestamp 1644511149
transform 1 0 81788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_889
timestamp 1644511149
transform 1 0 82892 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_895
timestamp 1644511149
transform 1 0 83444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_897
timestamp 1644511149
transform 1 0 83628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_909
timestamp 1644511149
transform 1 0 84732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_921
timestamp 1644511149
transform 1 0 85836 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_933
timestamp 1644511149
transform 1 0 86940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_945
timestamp 1644511149
transform 1 0 88044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_951
timestamp 1644511149
transform 1 0 88596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_953
timestamp 1644511149
transform 1 0 88780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_965
timestamp 1644511149
transform 1 0 89884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_977
timestamp 1644511149
transform 1 0 90988 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_989
timestamp 1644511149
transform 1 0 92092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1001
timestamp 1644511149
transform 1 0 93196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1007
timestamp 1644511149
transform 1 0 93748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1009
timestamp 1644511149
transform 1 0 93932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1021
timestamp 1644511149
transform 1 0 95036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1033
timestamp 1644511149
transform 1 0 96140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1045
timestamp 1644511149
transform 1 0 97244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1057
timestamp 1644511149
transform 1 0 98348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1063
timestamp 1644511149
transform 1 0 98900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1065
timestamp 1644511149
transform 1 0 99084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1077
timestamp 1644511149
transform 1 0 100188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1089
timestamp 1644511149
transform 1 0 101292 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1101
timestamp 1644511149
transform 1 0 102396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1113
timestamp 1644511149
transform 1 0 103500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1119
timestamp 1644511149
transform 1 0 104052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1121
timestamp 1644511149
transform 1 0 104236 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1133
timestamp 1644511149
transform 1 0 105340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1145
timestamp 1644511149
transform 1 0 106444 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1157
timestamp 1644511149
transform 1 0 107548 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1169
timestamp 1644511149
transform 1 0 108652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1175
timestamp 1644511149
transform 1 0 109204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1177
timestamp 1644511149
transform 1 0 109388 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1189
timestamp 1644511149
transform 1 0 110492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1201
timestamp 1644511149
transform 1 0 111596 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1213
timestamp 1644511149
transform 1 0 112700 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1225
timestamp 1644511149
transform 1 0 113804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1231
timestamp 1644511149
transform 1 0 114356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1233
timestamp 1644511149
transform 1 0 114540 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1245
timestamp 1644511149
transform 1 0 115644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1257
timestamp 1644511149
transform 1 0 116748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1269
timestamp 1644511149
transform 1 0 117852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1644511149
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1644511149
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1644511149
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1644511149
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_737
timestamp 1644511149
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1644511149
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1644511149
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_757
timestamp 1644511149
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_769
timestamp 1644511149
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_781
timestamp 1644511149
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_793
timestamp 1644511149
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1644511149
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1644511149
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_813
timestamp 1644511149
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_825
timestamp 1644511149
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_837
timestamp 1644511149
transform 1 0 78108 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_849
timestamp 1644511149
transform 1 0 79212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_861
timestamp 1644511149
transform 1 0 80316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_867
timestamp 1644511149
transform 1 0 80868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_869
timestamp 1644511149
transform 1 0 81052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_881
timestamp 1644511149
transform 1 0 82156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_893
timestamp 1644511149
transform 1 0 83260 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_905
timestamp 1644511149
transform 1 0 84364 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_917
timestamp 1644511149
transform 1 0 85468 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_923
timestamp 1644511149
transform 1 0 86020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_925
timestamp 1644511149
transform 1 0 86204 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_937
timestamp 1644511149
transform 1 0 87308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_949
timestamp 1644511149
transform 1 0 88412 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_961
timestamp 1644511149
transform 1 0 89516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_973
timestamp 1644511149
transform 1 0 90620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_979
timestamp 1644511149
transform 1 0 91172 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_981
timestamp 1644511149
transform 1 0 91356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_993
timestamp 1644511149
transform 1 0 92460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1005
timestamp 1644511149
transform 1 0 93564 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1017
timestamp 1644511149
transform 1 0 94668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1029
timestamp 1644511149
transform 1 0 95772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1035
timestamp 1644511149
transform 1 0 96324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1037
timestamp 1644511149
transform 1 0 96508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1049
timestamp 1644511149
transform 1 0 97612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1061
timestamp 1644511149
transform 1 0 98716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1073
timestamp 1644511149
transform 1 0 99820 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1085
timestamp 1644511149
transform 1 0 100924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1091
timestamp 1644511149
transform 1 0 101476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1093
timestamp 1644511149
transform 1 0 101660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1105
timestamp 1644511149
transform 1 0 102764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1117
timestamp 1644511149
transform 1 0 103868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1129
timestamp 1644511149
transform 1 0 104972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1141
timestamp 1644511149
transform 1 0 106076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1147
timestamp 1644511149
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1149
timestamp 1644511149
transform 1 0 106812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1161
timestamp 1644511149
transform 1 0 107916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1173
timestamp 1644511149
transform 1 0 109020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1185
timestamp 1644511149
transform 1 0 110124 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1197
timestamp 1644511149
transform 1 0 111228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1203
timestamp 1644511149
transform 1 0 111780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1205
timestamp 1644511149
transform 1 0 111964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1217
timestamp 1644511149
transform 1 0 113068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1229
timestamp 1644511149
transform 1 0 114172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1241
timestamp 1644511149
transform 1 0 115276 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1253
timestamp 1644511149
transform 1 0 116380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1259
timestamp 1644511149
transform 1 0 116932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1261
timestamp 1644511149
transform 1 0 117116 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_1273
timestamp 1644511149
transform 1 0 118220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1644511149
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1644511149
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_709
timestamp 1644511149
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1644511149
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1644511149
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_741
timestamp 1644511149
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_753
timestamp 1644511149
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_765
timestamp 1644511149
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1644511149
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1644511149
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_785
timestamp 1644511149
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_797
timestamp 1644511149
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_809
timestamp 1644511149
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_821
timestamp 1644511149
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1644511149
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1644511149
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_841
timestamp 1644511149
transform 1 0 78476 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_853
timestamp 1644511149
transform 1 0 79580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_865
timestamp 1644511149
transform 1 0 80684 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_877
timestamp 1644511149
transform 1 0 81788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_889
timestamp 1644511149
transform 1 0 82892 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_895
timestamp 1644511149
transform 1 0 83444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_897
timestamp 1644511149
transform 1 0 83628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_909
timestamp 1644511149
transform 1 0 84732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_921
timestamp 1644511149
transform 1 0 85836 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_933
timestamp 1644511149
transform 1 0 86940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_945
timestamp 1644511149
transform 1 0 88044 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_951
timestamp 1644511149
transform 1 0 88596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_953
timestamp 1644511149
transform 1 0 88780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_965
timestamp 1644511149
transform 1 0 89884 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_977
timestamp 1644511149
transform 1 0 90988 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_989
timestamp 1644511149
transform 1 0 92092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1001
timestamp 1644511149
transform 1 0 93196 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1007
timestamp 1644511149
transform 1 0 93748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1009
timestamp 1644511149
transform 1 0 93932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1021
timestamp 1644511149
transform 1 0 95036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1033
timestamp 1644511149
transform 1 0 96140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1045
timestamp 1644511149
transform 1 0 97244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1057
timestamp 1644511149
transform 1 0 98348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1063
timestamp 1644511149
transform 1 0 98900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1065
timestamp 1644511149
transform 1 0 99084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1077
timestamp 1644511149
transform 1 0 100188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1089
timestamp 1644511149
transform 1 0 101292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1101
timestamp 1644511149
transform 1 0 102396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1113
timestamp 1644511149
transform 1 0 103500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1119
timestamp 1644511149
transform 1 0 104052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1121
timestamp 1644511149
transform 1 0 104236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1133
timestamp 1644511149
transform 1 0 105340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1145
timestamp 1644511149
transform 1 0 106444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1157
timestamp 1644511149
transform 1 0 107548 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1169
timestamp 1644511149
transform 1 0 108652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1175
timestamp 1644511149
transform 1 0 109204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1177
timestamp 1644511149
transform 1 0 109388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1189
timestamp 1644511149
transform 1 0 110492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1201
timestamp 1644511149
transform 1 0 111596 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1213
timestamp 1644511149
transform 1 0 112700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1225
timestamp 1644511149
transform 1 0 113804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1231
timestamp 1644511149
transform 1 0 114356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1233
timestamp 1644511149
transform 1 0 114540 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1245
timestamp 1644511149
transform 1 0 115644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1257
timestamp 1644511149
transform 1 0 116748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1269
timestamp 1644511149
transform 1 0 117852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_625
timestamp 1644511149
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1644511149
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1644511149
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1644511149
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1644511149
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1644511149
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1644511149
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_725
timestamp 1644511149
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_737
timestamp 1644511149
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1644511149
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1644511149
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_757
timestamp 1644511149
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_769
timestamp 1644511149
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_781
timestamp 1644511149
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_793
timestamp 1644511149
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1644511149
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1644511149
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_813
timestamp 1644511149
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_825
timestamp 1644511149
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_837
timestamp 1644511149
transform 1 0 78108 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_849
timestamp 1644511149
transform 1 0 79212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_861
timestamp 1644511149
transform 1 0 80316 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_867
timestamp 1644511149
transform 1 0 80868 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_869
timestamp 1644511149
transform 1 0 81052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_881
timestamp 1644511149
transform 1 0 82156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_893
timestamp 1644511149
transform 1 0 83260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_905
timestamp 1644511149
transform 1 0 84364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_917
timestamp 1644511149
transform 1 0 85468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_923
timestamp 1644511149
transform 1 0 86020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_925
timestamp 1644511149
transform 1 0 86204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_937
timestamp 1644511149
transform 1 0 87308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_949
timestamp 1644511149
transform 1 0 88412 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_961
timestamp 1644511149
transform 1 0 89516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_973
timestamp 1644511149
transform 1 0 90620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_979
timestamp 1644511149
transform 1 0 91172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_981
timestamp 1644511149
transform 1 0 91356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_993
timestamp 1644511149
transform 1 0 92460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1005
timestamp 1644511149
transform 1 0 93564 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1017
timestamp 1644511149
transform 1 0 94668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1029
timestamp 1644511149
transform 1 0 95772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1035
timestamp 1644511149
transform 1 0 96324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1037
timestamp 1644511149
transform 1 0 96508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1049
timestamp 1644511149
transform 1 0 97612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1061
timestamp 1644511149
transform 1 0 98716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1073
timestamp 1644511149
transform 1 0 99820 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1085
timestamp 1644511149
transform 1 0 100924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1091
timestamp 1644511149
transform 1 0 101476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1093
timestamp 1644511149
transform 1 0 101660 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1105
timestamp 1644511149
transform 1 0 102764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1117
timestamp 1644511149
transform 1 0 103868 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1129
timestamp 1644511149
transform 1 0 104972 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1141
timestamp 1644511149
transform 1 0 106076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1147
timestamp 1644511149
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1149
timestamp 1644511149
transform 1 0 106812 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1161
timestamp 1644511149
transform 1 0 107916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1173
timestamp 1644511149
transform 1 0 109020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1185
timestamp 1644511149
transform 1 0 110124 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1197
timestamp 1644511149
transform 1 0 111228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1203
timestamp 1644511149
transform 1 0 111780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1205
timestamp 1644511149
transform 1 0 111964 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1217
timestamp 1644511149
transform 1 0 113068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1229
timestamp 1644511149
transform 1 0 114172 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1241
timestamp 1644511149
transform 1 0 115276 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1253
timestamp 1644511149
transform 1 0 116380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1259
timestamp 1644511149
transform 1 0 116932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1261
timestamp 1644511149
transform 1 0 117116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_1273
timestamp 1644511149
transform 1 0 118220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_9
timestamp 1644511149
transform 1 0 1932 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_21
timestamp 1644511149
transform 1 0 3036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_33
timestamp 1644511149
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1644511149
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1644511149
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_741
timestamp 1644511149
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_753
timestamp 1644511149
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_765
timestamp 1644511149
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1644511149
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1644511149
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_785
timestamp 1644511149
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_797
timestamp 1644511149
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_809
timestamp 1644511149
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_821
timestamp 1644511149
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1644511149
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1644511149
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_841
timestamp 1644511149
transform 1 0 78476 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_853
timestamp 1644511149
transform 1 0 79580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_865
timestamp 1644511149
transform 1 0 80684 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_877
timestamp 1644511149
transform 1 0 81788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_889
timestamp 1644511149
transform 1 0 82892 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_895
timestamp 1644511149
transform 1 0 83444 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_897
timestamp 1644511149
transform 1 0 83628 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_909
timestamp 1644511149
transform 1 0 84732 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_921
timestamp 1644511149
transform 1 0 85836 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_933
timestamp 1644511149
transform 1 0 86940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_945
timestamp 1644511149
transform 1 0 88044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_951
timestamp 1644511149
transform 1 0 88596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_953
timestamp 1644511149
transform 1 0 88780 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_965
timestamp 1644511149
transform 1 0 89884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_977
timestamp 1644511149
transform 1 0 90988 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_989
timestamp 1644511149
transform 1 0 92092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1001
timestamp 1644511149
transform 1 0 93196 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1007
timestamp 1644511149
transform 1 0 93748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1009
timestamp 1644511149
transform 1 0 93932 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1021
timestamp 1644511149
transform 1 0 95036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1033
timestamp 1644511149
transform 1 0 96140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1045
timestamp 1644511149
transform 1 0 97244 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1057
timestamp 1644511149
transform 1 0 98348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1063
timestamp 1644511149
transform 1 0 98900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1065
timestamp 1644511149
transform 1 0 99084 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1077
timestamp 1644511149
transform 1 0 100188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1089
timestamp 1644511149
transform 1 0 101292 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1101
timestamp 1644511149
transform 1 0 102396 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1113
timestamp 1644511149
transform 1 0 103500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1119
timestamp 1644511149
transform 1 0 104052 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1121
timestamp 1644511149
transform 1 0 104236 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1133
timestamp 1644511149
transform 1 0 105340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1145
timestamp 1644511149
transform 1 0 106444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1157
timestamp 1644511149
transform 1 0 107548 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1169
timestamp 1644511149
transform 1 0 108652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1175
timestamp 1644511149
transform 1 0 109204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1177
timestamp 1644511149
transform 1 0 109388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1189
timestamp 1644511149
transform 1 0 110492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1201
timestamp 1644511149
transform 1 0 111596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1213
timestamp 1644511149
transform 1 0 112700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1225
timestamp 1644511149
transform 1 0 113804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1231
timestamp 1644511149
transform 1 0 114356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1233
timestamp 1644511149
transform 1 0 114540 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1245
timestamp 1644511149
transform 1 0 115644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1257
timestamp 1644511149
transform 1 0 116748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1267
timestamp 1644511149
transform 1 0 117668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_1273
timestamp 1644511149
transform 1 0 118220 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_713
timestamp 1644511149
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_725
timestamp 1644511149
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_737
timestamp 1644511149
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1644511149
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1644511149
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_757
timestamp 1644511149
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_769
timestamp 1644511149
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_781
timestamp 1644511149
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_793
timestamp 1644511149
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1644511149
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1644511149
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_813
timestamp 1644511149
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_825
timestamp 1644511149
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_837
timestamp 1644511149
transform 1 0 78108 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_849
timestamp 1644511149
transform 1 0 79212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_861
timestamp 1644511149
transform 1 0 80316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_867
timestamp 1644511149
transform 1 0 80868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_869
timestamp 1644511149
transform 1 0 81052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_881
timestamp 1644511149
transform 1 0 82156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_893
timestamp 1644511149
transform 1 0 83260 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_905
timestamp 1644511149
transform 1 0 84364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_917
timestamp 1644511149
transform 1 0 85468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_923
timestamp 1644511149
transform 1 0 86020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_925
timestamp 1644511149
transform 1 0 86204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_937
timestamp 1644511149
transform 1 0 87308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_949
timestamp 1644511149
transform 1 0 88412 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_961
timestamp 1644511149
transform 1 0 89516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_973
timestamp 1644511149
transform 1 0 90620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_979
timestamp 1644511149
transform 1 0 91172 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_981
timestamp 1644511149
transform 1 0 91356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_993
timestamp 1644511149
transform 1 0 92460 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1005
timestamp 1644511149
transform 1 0 93564 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1017
timestamp 1644511149
transform 1 0 94668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1029
timestamp 1644511149
transform 1 0 95772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1035
timestamp 1644511149
transform 1 0 96324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1037
timestamp 1644511149
transform 1 0 96508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1049
timestamp 1644511149
transform 1 0 97612 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1061
timestamp 1644511149
transform 1 0 98716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1073
timestamp 1644511149
transform 1 0 99820 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1085
timestamp 1644511149
transform 1 0 100924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1091
timestamp 1644511149
transform 1 0 101476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1093
timestamp 1644511149
transform 1 0 101660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1105
timestamp 1644511149
transform 1 0 102764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1117
timestamp 1644511149
transform 1 0 103868 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1129
timestamp 1644511149
transform 1 0 104972 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1141
timestamp 1644511149
transform 1 0 106076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1147
timestamp 1644511149
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1149
timestamp 1644511149
transform 1 0 106812 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1161
timestamp 1644511149
transform 1 0 107916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1173
timestamp 1644511149
transform 1 0 109020 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1185
timestamp 1644511149
transform 1 0 110124 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1197
timestamp 1644511149
transform 1 0 111228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1203
timestamp 1644511149
transform 1 0 111780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1205
timestamp 1644511149
transform 1 0 111964 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1217
timestamp 1644511149
transform 1 0 113068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1229
timestamp 1644511149
transform 1 0 114172 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1241
timestamp 1644511149
transform 1 0 115276 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1253
timestamp 1644511149
transform 1 0 116380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1259
timestamp 1644511149
transform 1 0 116932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1261
timestamp 1644511149
transform 1 0 117116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_1273
timestamp 1644511149
transform 1 0 118220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1644511149
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_741
timestamp 1644511149
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_753
timestamp 1644511149
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_765
timestamp 1644511149
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1644511149
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1644511149
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_785
timestamp 1644511149
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_797
timestamp 1644511149
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_809
timestamp 1644511149
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_821
timestamp 1644511149
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1644511149
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1644511149
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_841
timestamp 1644511149
transform 1 0 78476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_853
timestamp 1644511149
transform 1 0 79580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_865
timestamp 1644511149
transform 1 0 80684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_877
timestamp 1644511149
transform 1 0 81788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_889
timestamp 1644511149
transform 1 0 82892 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_895
timestamp 1644511149
transform 1 0 83444 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_897
timestamp 1644511149
transform 1 0 83628 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_909
timestamp 1644511149
transform 1 0 84732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_921
timestamp 1644511149
transform 1 0 85836 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_933
timestamp 1644511149
transform 1 0 86940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_945
timestamp 1644511149
transform 1 0 88044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_951
timestamp 1644511149
transform 1 0 88596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_953
timestamp 1644511149
transform 1 0 88780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_965
timestamp 1644511149
transform 1 0 89884 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_977
timestamp 1644511149
transform 1 0 90988 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_989
timestamp 1644511149
transform 1 0 92092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1001
timestamp 1644511149
transform 1 0 93196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1007
timestamp 1644511149
transform 1 0 93748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1009
timestamp 1644511149
transform 1 0 93932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1021
timestamp 1644511149
transform 1 0 95036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1033
timestamp 1644511149
transform 1 0 96140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1045
timestamp 1644511149
transform 1 0 97244 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1057
timestamp 1644511149
transform 1 0 98348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1063
timestamp 1644511149
transform 1 0 98900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1065
timestamp 1644511149
transform 1 0 99084 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1077
timestamp 1644511149
transform 1 0 100188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1089
timestamp 1644511149
transform 1 0 101292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1101
timestamp 1644511149
transform 1 0 102396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1113
timestamp 1644511149
transform 1 0 103500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1119
timestamp 1644511149
transform 1 0 104052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1121
timestamp 1644511149
transform 1 0 104236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1133
timestamp 1644511149
transform 1 0 105340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1145
timestamp 1644511149
transform 1 0 106444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1157
timestamp 1644511149
transform 1 0 107548 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1169
timestamp 1644511149
transform 1 0 108652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1175
timestamp 1644511149
transform 1 0 109204 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1177
timestamp 1644511149
transform 1 0 109388 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1189
timestamp 1644511149
transform 1 0 110492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1201
timestamp 1644511149
transform 1 0 111596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1213
timestamp 1644511149
transform 1 0 112700 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1225
timestamp 1644511149
transform 1 0 113804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1231
timestamp 1644511149
transform 1 0 114356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1233
timestamp 1644511149
transform 1 0 114540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1245
timestamp 1644511149
transform 1 0 115644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1257
timestamp 1644511149
transform 1 0 116748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_1267
timestamp 1644511149
transform 1 0 117668 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1273
timestamp 1644511149
transform 1 0 118220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1644511149
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_737
timestamp 1644511149
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1644511149
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1644511149
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_757
timestamp 1644511149
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_769
timestamp 1644511149
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_781
timestamp 1644511149
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_793
timestamp 1644511149
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1644511149
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1644511149
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_813
timestamp 1644511149
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_825
timestamp 1644511149
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_837
timestamp 1644511149
transform 1 0 78108 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_849
timestamp 1644511149
transform 1 0 79212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_861
timestamp 1644511149
transform 1 0 80316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_867
timestamp 1644511149
transform 1 0 80868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_869
timestamp 1644511149
transform 1 0 81052 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_881
timestamp 1644511149
transform 1 0 82156 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_893
timestamp 1644511149
transform 1 0 83260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_905
timestamp 1644511149
transform 1 0 84364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_917
timestamp 1644511149
transform 1 0 85468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_923
timestamp 1644511149
transform 1 0 86020 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_925
timestamp 1644511149
transform 1 0 86204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_937
timestamp 1644511149
transform 1 0 87308 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_949
timestamp 1644511149
transform 1 0 88412 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_961
timestamp 1644511149
transform 1 0 89516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_973
timestamp 1644511149
transform 1 0 90620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_979
timestamp 1644511149
transform 1 0 91172 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_981
timestamp 1644511149
transform 1 0 91356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_993
timestamp 1644511149
transform 1 0 92460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1005
timestamp 1644511149
transform 1 0 93564 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1017
timestamp 1644511149
transform 1 0 94668 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1029
timestamp 1644511149
transform 1 0 95772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1035
timestamp 1644511149
transform 1 0 96324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1037
timestamp 1644511149
transform 1 0 96508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1049
timestamp 1644511149
transform 1 0 97612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1061
timestamp 1644511149
transform 1 0 98716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1073
timestamp 1644511149
transform 1 0 99820 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1085
timestamp 1644511149
transform 1 0 100924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1091
timestamp 1644511149
transform 1 0 101476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1093
timestamp 1644511149
transform 1 0 101660 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1105
timestamp 1644511149
transform 1 0 102764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1117
timestamp 1644511149
transform 1 0 103868 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1129
timestamp 1644511149
transform 1 0 104972 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1141
timestamp 1644511149
transform 1 0 106076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1147
timestamp 1644511149
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1149
timestamp 1644511149
transform 1 0 106812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1161
timestamp 1644511149
transform 1 0 107916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1173
timestamp 1644511149
transform 1 0 109020 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1185
timestamp 1644511149
transform 1 0 110124 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1197
timestamp 1644511149
transform 1 0 111228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1203
timestamp 1644511149
transform 1 0 111780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1205
timestamp 1644511149
transform 1 0 111964 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1217
timestamp 1644511149
transform 1 0 113068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1229
timestamp 1644511149
transform 1 0 114172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1241
timestamp 1644511149
transform 1 0 115276 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1253
timestamp 1644511149
transform 1 0 116380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1259
timestamp 1644511149
transform 1 0 116932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1261
timestamp 1644511149
transform 1 0 117116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_1273
timestamp 1644511149
transform 1 0 118220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_741
timestamp 1644511149
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_753
timestamp 1644511149
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_765
timestamp 1644511149
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1644511149
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1644511149
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_785
timestamp 1644511149
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_797
timestamp 1644511149
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_809
timestamp 1644511149
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_821
timestamp 1644511149
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_833
timestamp 1644511149
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_839
timestamp 1644511149
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_841
timestamp 1644511149
transform 1 0 78476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_853
timestamp 1644511149
transform 1 0 79580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_865
timestamp 1644511149
transform 1 0 80684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_877
timestamp 1644511149
transform 1 0 81788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_889
timestamp 1644511149
transform 1 0 82892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_895
timestamp 1644511149
transform 1 0 83444 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_897
timestamp 1644511149
transform 1 0 83628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_909
timestamp 1644511149
transform 1 0 84732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_921
timestamp 1644511149
transform 1 0 85836 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_933
timestamp 1644511149
transform 1 0 86940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_945
timestamp 1644511149
transform 1 0 88044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_951
timestamp 1644511149
transform 1 0 88596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_953
timestamp 1644511149
transform 1 0 88780 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_965
timestamp 1644511149
transform 1 0 89884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_977
timestamp 1644511149
transform 1 0 90988 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_989
timestamp 1644511149
transform 1 0 92092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1001
timestamp 1644511149
transform 1 0 93196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1007
timestamp 1644511149
transform 1 0 93748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1009
timestamp 1644511149
transform 1 0 93932 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1021
timestamp 1644511149
transform 1 0 95036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1033
timestamp 1644511149
transform 1 0 96140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1045
timestamp 1644511149
transform 1 0 97244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1057
timestamp 1644511149
transform 1 0 98348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1063
timestamp 1644511149
transform 1 0 98900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1065
timestamp 1644511149
transform 1 0 99084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1077
timestamp 1644511149
transform 1 0 100188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1089
timestamp 1644511149
transform 1 0 101292 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1101
timestamp 1644511149
transform 1 0 102396 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1113
timestamp 1644511149
transform 1 0 103500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1119
timestamp 1644511149
transform 1 0 104052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1121
timestamp 1644511149
transform 1 0 104236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1133
timestamp 1644511149
transform 1 0 105340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1145
timestamp 1644511149
transform 1 0 106444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1157
timestamp 1644511149
transform 1 0 107548 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1169
timestamp 1644511149
transform 1 0 108652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1175
timestamp 1644511149
transform 1 0 109204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1177
timestamp 1644511149
transform 1 0 109388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1189
timestamp 1644511149
transform 1 0 110492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1201
timestamp 1644511149
transform 1 0 111596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1213
timestamp 1644511149
transform 1 0 112700 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1225
timestamp 1644511149
transform 1 0 113804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1231
timestamp 1644511149
transform 1 0 114356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1233
timestamp 1644511149
transform 1 0 114540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1245
timestamp 1644511149
transform 1 0 115644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1257
timestamp 1644511149
transform 1 0 116748 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1269
timestamp 1644511149
transform 1 0 117852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_737
timestamp 1644511149
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1644511149
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1644511149
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_757
timestamp 1644511149
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_769
timestamp 1644511149
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_781
timestamp 1644511149
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_793
timestamp 1644511149
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1644511149
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1644511149
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_813
timestamp 1644511149
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_825
timestamp 1644511149
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_837
timestamp 1644511149
transform 1 0 78108 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_849
timestamp 1644511149
transform 1 0 79212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_861
timestamp 1644511149
transform 1 0 80316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_867
timestamp 1644511149
transform 1 0 80868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_869
timestamp 1644511149
transform 1 0 81052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_881
timestamp 1644511149
transform 1 0 82156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_893
timestamp 1644511149
transform 1 0 83260 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_905
timestamp 1644511149
transform 1 0 84364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_917
timestamp 1644511149
transform 1 0 85468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_923
timestamp 1644511149
transform 1 0 86020 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_925
timestamp 1644511149
transform 1 0 86204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_937
timestamp 1644511149
transform 1 0 87308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_949
timestamp 1644511149
transform 1 0 88412 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_961
timestamp 1644511149
transform 1 0 89516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_973
timestamp 1644511149
transform 1 0 90620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_979
timestamp 1644511149
transform 1 0 91172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_981
timestamp 1644511149
transform 1 0 91356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_993
timestamp 1644511149
transform 1 0 92460 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1005
timestamp 1644511149
transform 1 0 93564 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1017
timestamp 1644511149
transform 1 0 94668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1029
timestamp 1644511149
transform 1 0 95772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1035
timestamp 1644511149
transform 1 0 96324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1037
timestamp 1644511149
transform 1 0 96508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1049
timestamp 1644511149
transform 1 0 97612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1061
timestamp 1644511149
transform 1 0 98716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1073
timestamp 1644511149
transform 1 0 99820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1085
timestamp 1644511149
transform 1 0 100924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1091
timestamp 1644511149
transform 1 0 101476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1093
timestamp 1644511149
transform 1 0 101660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1105
timestamp 1644511149
transform 1 0 102764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1117
timestamp 1644511149
transform 1 0 103868 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1129
timestamp 1644511149
transform 1 0 104972 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1141
timestamp 1644511149
transform 1 0 106076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1147
timestamp 1644511149
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1149
timestamp 1644511149
transform 1 0 106812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1161
timestamp 1644511149
transform 1 0 107916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1173
timestamp 1644511149
transform 1 0 109020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1185
timestamp 1644511149
transform 1 0 110124 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1197
timestamp 1644511149
transform 1 0 111228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1203
timestamp 1644511149
transform 1 0 111780 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1205
timestamp 1644511149
transform 1 0 111964 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1217
timestamp 1644511149
transform 1 0 113068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1229
timestamp 1644511149
transform 1 0 114172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1241
timestamp 1644511149
transform 1 0 115276 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1253
timestamp 1644511149
transform 1 0 116380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1259
timestamp 1644511149
transform 1 0 116932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1261
timestamp 1644511149
transform 1 0 117116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_1273
timestamp 1644511149
transform 1 0 118220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_9
timestamp 1644511149
transform 1 0 1932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_21
timestamp 1644511149
transform 1 0 3036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_33
timestamp 1644511149
transform 1 0 4140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_45
timestamp 1644511149
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1644511149
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_629
timestamp 1644511149
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_641
timestamp 1644511149
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_653
timestamp 1644511149
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1644511149
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_741
timestamp 1644511149
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_753
timestamp 1644511149
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_765
timestamp 1644511149
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1644511149
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1644511149
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_785
timestamp 1644511149
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_797
timestamp 1644511149
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_809
timestamp 1644511149
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_821
timestamp 1644511149
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_833
timestamp 1644511149
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_839
timestamp 1644511149
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_841
timestamp 1644511149
transform 1 0 78476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_853
timestamp 1644511149
transform 1 0 79580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_865
timestamp 1644511149
transform 1 0 80684 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_877
timestamp 1644511149
transform 1 0 81788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_889
timestamp 1644511149
transform 1 0 82892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_895
timestamp 1644511149
transform 1 0 83444 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_897
timestamp 1644511149
transform 1 0 83628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_909
timestamp 1644511149
transform 1 0 84732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_921
timestamp 1644511149
transform 1 0 85836 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_933
timestamp 1644511149
transform 1 0 86940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_945
timestamp 1644511149
transform 1 0 88044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_951
timestamp 1644511149
transform 1 0 88596 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_953
timestamp 1644511149
transform 1 0 88780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_965
timestamp 1644511149
transform 1 0 89884 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_977
timestamp 1644511149
transform 1 0 90988 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_989
timestamp 1644511149
transform 1 0 92092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1001
timestamp 1644511149
transform 1 0 93196 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1007
timestamp 1644511149
transform 1 0 93748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1009
timestamp 1644511149
transform 1 0 93932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1021
timestamp 1644511149
transform 1 0 95036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1033
timestamp 1644511149
transform 1 0 96140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1045
timestamp 1644511149
transform 1 0 97244 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1057
timestamp 1644511149
transform 1 0 98348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1063
timestamp 1644511149
transform 1 0 98900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1065
timestamp 1644511149
transform 1 0 99084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1077
timestamp 1644511149
transform 1 0 100188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1089
timestamp 1644511149
transform 1 0 101292 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1101
timestamp 1644511149
transform 1 0 102396 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1113
timestamp 1644511149
transform 1 0 103500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1119
timestamp 1644511149
transform 1 0 104052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1121
timestamp 1644511149
transform 1 0 104236 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1133
timestamp 1644511149
transform 1 0 105340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1145
timestamp 1644511149
transform 1 0 106444 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1157
timestamp 1644511149
transform 1 0 107548 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1169
timestamp 1644511149
transform 1 0 108652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1175
timestamp 1644511149
transform 1 0 109204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1177
timestamp 1644511149
transform 1 0 109388 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1189
timestamp 1644511149
transform 1 0 110492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1201
timestamp 1644511149
transform 1 0 111596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1213
timestamp 1644511149
transform 1 0 112700 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1225
timestamp 1644511149
transform 1 0 113804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1231
timestamp 1644511149
transform 1 0 114356 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1233
timestamp 1644511149
transform 1 0 114540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1245
timestamp 1644511149
transform 1 0 115644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1257
timestamp 1644511149
transform 1 0 116748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1269
timestamp 1644511149
transform 1 0 117852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_625
timestamp 1644511149
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1644511149
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1644511149
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_737
timestamp 1644511149
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1644511149
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1644511149
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_757
timestamp 1644511149
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_769
timestamp 1644511149
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_781
timestamp 1644511149
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_793
timestamp 1644511149
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1644511149
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1644511149
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_813
timestamp 1644511149
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_825
timestamp 1644511149
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_837
timestamp 1644511149
transform 1 0 78108 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_849
timestamp 1644511149
transform 1 0 79212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_861
timestamp 1644511149
transform 1 0 80316 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_867
timestamp 1644511149
transform 1 0 80868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_869
timestamp 1644511149
transform 1 0 81052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_881
timestamp 1644511149
transform 1 0 82156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_893
timestamp 1644511149
transform 1 0 83260 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_905
timestamp 1644511149
transform 1 0 84364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_917
timestamp 1644511149
transform 1 0 85468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_923
timestamp 1644511149
transform 1 0 86020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_925
timestamp 1644511149
transform 1 0 86204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_937
timestamp 1644511149
transform 1 0 87308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_949
timestamp 1644511149
transform 1 0 88412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_961
timestamp 1644511149
transform 1 0 89516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_973
timestamp 1644511149
transform 1 0 90620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_979
timestamp 1644511149
transform 1 0 91172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_981
timestamp 1644511149
transform 1 0 91356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_993
timestamp 1644511149
transform 1 0 92460 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1005
timestamp 1644511149
transform 1 0 93564 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1017
timestamp 1644511149
transform 1 0 94668 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1029
timestamp 1644511149
transform 1 0 95772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1035
timestamp 1644511149
transform 1 0 96324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1037
timestamp 1644511149
transform 1 0 96508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1049
timestamp 1644511149
transform 1 0 97612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1061
timestamp 1644511149
transform 1 0 98716 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1073
timestamp 1644511149
transform 1 0 99820 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1085
timestamp 1644511149
transform 1 0 100924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1091
timestamp 1644511149
transform 1 0 101476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1093
timestamp 1644511149
transform 1 0 101660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1105
timestamp 1644511149
transform 1 0 102764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1117
timestamp 1644511149
transform 1 0 103868 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1129
timestamp 1644511149
transform 1 0 104972 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1141
timestamp 1644511149
transform 1 0 106076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1147
timestamp 1644511149
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1149
timestamp 1644511149
transform 1 0 106812 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1161
timestamp 1644511149
transform 1 0 107916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1173
timestamp 1644511149
transform 1 0 109020 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1185
timestamp 1644511149
transform 1 0 110124 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1197
timestamp 1644511149
transform 1 0 111228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1203
timestamp 1644511149
transform 1 0 111780 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1205
timestamp 1644511149
transform 1 0 111964 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1217
timestamp 1644511149
transform 1 0 113068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1229
timestamp 1644511149
transform 1 0 114172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1241
timestamp 1644511149
transform 1 0 115276 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1253
timestamp 1644511149
transform 1 0 116380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1259
timestamp 1644511149
transform 1 0 116932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1261
timestamp 1644511149
transform 1 0 117116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_1273
timestamp 1644511149
transform 1 0 118220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_629
timestamp 1644511149
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_641
timestamp 1644511149
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_653
timestamp 1644511149
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1644511149
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1644511149
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_741
timestamp 1644511149
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_753
timestamp 1644511149
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_765
timestamp 1644511149
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1644511149
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1644511149
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_785
timestamp 1644511149
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_797
timestamp 1644511149
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_809
timestamp 1644511149
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_821
timestamp 1644511149
transform 1 0 76636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_833
timestamp 1644511149
transform 1 0 77740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_839
timestamp 1644511149
transform 1 0 78292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_841
timestamp 1644511149
transform 1 0 78476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_853
timestamp 1644511149
transform 1 0 79580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_865
timestamp 1644511149
transform 1 0 80684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_877
timestamp 1644511149
transform 1 0 81788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_889
timestamp 1644511149
transform 1 0 82892 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_895
timestamp 1644511149
transform 1 0 83444 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_897
timestamp 1644511149
transform 1 0 83628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_909
timestamp 1644511149
transform 1 0 84732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_921
timestamp 1644511149
transform 1 0 85836 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_933
timestamp 1644511149
transform 1 0 86940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_945
timestamp 1644511149
transform 1 0 88044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_951
timestamp 1644511149
transform 1 0 88596 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_953
timestamp 1644511149
transform 1 0 88780 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_965
timestamp 1644511149
transform 1 0 89884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_977
timestamp 1644511149
transform 1 0 90988 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_989
timestamp 1644511149
transform 1 0 92092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1001
timestamp 1644511149
transform 1 0 93196 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1007
timestamp 1644511149
transform 1 0 93748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1009
timestamp 1644511149
transform 1 0 93932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1021
timestamp 1644511149
transform 1 0 95036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1033
timestamp 1644511149
transform 1 0 96140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1045
timestamp 1644511149
transform 1 0 97244 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1057
timestamp 1644511149
transform 1 0 98348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1063
timestamp 1644511149
transform 1 0 98900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1065
timestamp 1644511149
transform 1 0 99084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1077
timestamp 1644511149
transform 1 0 100188 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1089
timestamp 1644511149
transform 1 0 101292 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1101
timestamp 1644511149
transform 1 0 102396 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1113
timestamp 1644511149
transform 1 0 103500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1119
timestamp 1644511149
transform 1 0 104052 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1121
timestamp 1644511149
transform 1 0 104236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1133
timestamp 1644511149
transform 1 0 105340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1145
timestamp 1644511149
transform 1 0 106444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1157
timestamp 1644511149
transform 1 0 107548 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1169
timestamp 1644511149
transform 1 0 108652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1175
timestamp 1644511149
transform 1 0 109204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1177
timestamp 1644511149
transform 1 0 109388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1189
timestamp 1644511149
transform 1 0 110492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1201
timestamp 1644511149
transform 1 0 111596 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1213
timestamp 1644511149
transform 1 0 112700 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1225
timestamp 1644511149
transform 1 0 113804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1231
timestamp 1644511149
transform 1 0 114356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1233
timestamp 1644511149
transform 1 0 114540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1245
timestamp 1644511149
transform 1 0 115644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_1257
timestamp 1644511149
transform 1 0 116748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_1267
timestamp 1644511149
transform 1 0 117668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1273
timestamp 1644511149
transform 1 0 118220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_625
timestamp 1644511149
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1644511149
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1644511149
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1644511149
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1644511149
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1644511149
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1644511149
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_737
timestamp 1644511149
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1644511149
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1644511149
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_757
timestamp 1644511149
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_769
timestamp 1644511149
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_781
timestamp 1644511149
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_793
timestamp 1644511149
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1644511149
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1644511149
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_813
timestamp 1644511149
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_825
timestamp 1644511149
transform 1 0 77004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_837
timestamp 1644511149
transform 1 0 78108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_849
timestamp 1644511149
transform 1 0 79212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_861
timestamp 1644511149
transform 1 0 80316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_867
timestamp 1644511149
transform 1 0 80868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_869
timestamp 1644511149
transform 1 0 81052 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_881
timestamp 1644511149
transform 1 0 82156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_893
timestamp 1644511149
transform 1 0 83260 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_905
timestamp 1644511149
transform 1 0 84364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_917
timestamp 1644511149
transform 1 0 85468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_923
timestamp 1644511149
transform 1 0 86020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_925
timestamp 1644511149
transform 1 0 86204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_937
timestamp 1644511149
transform 1 0 87308 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_949
timestamp 1644511149
transform 1 0 88412 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_961
timestamp 1644511149
transform 1 0 89516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_973
timestamp 1644511149
transform 1 0 90620 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_979
timestamp 1644511149
transform 1 0 91172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_981
timestamp 1644511149
transform 1 0 91356 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_993
timestamp 1644511149
transform 1 0 92460 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1005
timestamp 1644511149
transform 1 0 93564 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1017
timestamp 1644511149
transform 1 0 94668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1029
timestamp 1644511149
transform 1 0 95772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1035
timestamp 1644511149
transform 1 0 96324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1037
timestamp 1644511149
transform 1 0 96508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1049
timestamp 1644511149
transform 1 0 97612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1061
timestamp 1644511149
transform 1 0 98716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1073
timestamp 1644511149
transform 1 0 99820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1085
timestamp 1644511149
transform 1 0 100924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1091
timestamp 1644511149
transform 1 0 101476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1093
timestamp 1644511149
transform 1 0 101660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1105
timestamp 1644511149
transform 1 0 102764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1117
timestamp 1644511149
transform 1 0 103868 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1129
timestamp 1644511149
transform 1 0 104972 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1141
timestamp 1644511149
transform 1 0 106076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1147
timestamp 1644511149
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1149
timestamp 1644511149
transform 1 0 106812 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1161
timestamp 1644511149
transform 1 0 107916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1173
timestamp 1644511149
transform 1 0 109020 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1185
timestamp 1644511149
transform 1 0 110124 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1197
timestamp 1644511149
transform 1 0 111228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1203
timestamp 1644511149
transform 1 0 111780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1205
timestamp 1644511149
transform 1 0 111964 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1217
timestamp 1644511149
transform 1 0 113068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1229
timestamp 1644511149
transform 1 0 114172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1241
timestamp 1644511149
transform 1 0 115276 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1253
timestamp 1644511149
transform 1 0 116380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1259
timestamp 1644511149
transform 1 0 116932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1261
timestamp 1644511149
transform 1 0 117116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1273
timestamp 1644511149
transform 1 0 118220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_653
timestamp 1644511149
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1644511149
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1644511149
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_741
timestamp 1644511149
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_753
timestamp 1644511149
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_765
timestamp 1644511149
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1644511149
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1644511149
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_785
timestamp 1644511149
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_797
timestamp 1644511149
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_809
timestamp 1644511149
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_821
timestamp 1644511149
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_833
timestamp 1644511149
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_839
timestamp 1644511149
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_841
timestamp 1644511149
transform 1 0 78476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_853
timestamp 1644511149
transform 1 0 79580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_865
timestamp 1644511149
transform 1 0 80684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_877
timestamp 1644511149
transform 1 0 81788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_889
timestamp 1644511149
transform 1 0 82892 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_895
timestamp 1644511149
transform 1 0 83444 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_897
timestamp 1644511149
transform 1 0 83628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_909
timestamp 1644511149
transform 1 0 84732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_921
timestamp 1644511149
transform 1 0 85836 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_933
timestamp 1644511149
transform 1 0 86940 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_945
timestamp 1644511149
transform 1 0 88044 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_951
timestamp 1644511149
transform 1 0 88596 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_953
timestamp 1644511149
transform 1 0 88780 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_965
timestamp 1644511149
transform 1 0 89884 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_977
timestamp 1644511149
transform 1 0 90988 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_989
timestamp 1644511149
transform 1 0 92092 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1001
timestamp 1644511149
transform 1 0 93196 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1007
timestamp 1644511149
transform 1 0 93748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1009
timestamp 1644511149
transform 1 0 93932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1021
timestamp 1644511149
transform 1 0 95036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1033
timestamp 1644511149
transform 1 0 96140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1045
timestamp 1644511149
transform 1 0 97244 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1057
timestamp 1644511149
transform 1 0 98348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1063
timestamp 1644511149
transform 1 0 98900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1065
timestamp 1644511149
transform 1 0 99084 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1077
timestamp 1644511149
transform 1 0 100188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1089
timestamp 1644511149
transform 1 0 101292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1101
timestamp 1644511149
transform 1 0 102396 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1113
timestamp 1644511149
transform 1 0 103500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1119
timestamp 1644511149
transform 1 0 104052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1121
timestamp 1644511149
transform 1 0 104236 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1133
timestamp 1644511149
transform 1 0 105340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1145
timestamp 1644511149
transform 1 0 106444 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1157
timestamp 1644511149
transform 1 0 107548 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1169
timestamp 1644511149
transform 1 0 108652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1175
timestamp 1644511149
transform 1 0 109204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1177
timestamp 1644511149
transform 1 0 109388 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1189
timestamp 1644511149
transform 1 0 110492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1201
timestamp 1644511149
transform 1 0 111596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1213
timestamp 1644511149
transform 1 0 112700 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1225
timestamp 1644511149
transform 1 0 113804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1231
timestamp 1644511149
transform 1 0 114356 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1233
timestamp 1644511149
transform 1 0 114540 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1245
timestamp 1644511149
transform 1 0 115644 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1257
timestamp 1644511149
transform 1 0 116748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1269
timestamp 1644511149
transform 1 0 117852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1644511149
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1644511149
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1644511149
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1644511149
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1644511149
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_737
timestamp 1644511149
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1644511149
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1644511149
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_757
timestamp 1644511149
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_769
timestamp 1644511149
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_781
timestamp 1644511149
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_793
timestamp 1644511149
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1644511149
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1644511149
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_813
timestamp 1644511149
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_825
timestamp 1644511149
transform 1 0 77004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_837
timestamp 1644511149
transform 1 0 78108 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_849
timestamp 1644511149
transform 1 0 79212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_861
timestamp 1644511149
transform 1 0 80316 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_867
timestamp 1644511149
transform 1 0 80868 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_869
timestamp 1644511149
transform 1 0 81052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_881
timestamp 1644511149
transform 1 0 82156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_893
timestamp 1644511149
transform 1 0 83260 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_905
timestamp 1644511149
transform 1 0 84364 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_917
timestamp 1644511149
transform 1 0 85468 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_923
timestamp 1644511149
transform 1 0 86020 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_925
timestamp 1644511149
transform 1 0 86204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_937
timestamp 1644511149
transform 1 0 87308 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_949
timestamp 1644511149
transform 1 0 88412 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_961
timestamp 1644511149
transform 1 0 89516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_973
timestamp 1644511149
transform 1 0 90620 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_979
timestamp 1644511149
transform 1 0 91172 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_981
timestamp 1644511149
transform 1 0 91356 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_993
timestamp 1644511149
transform 1 0 92460 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1005
timestamp 1644511149
transform 1 0 93564 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1017
timestamp 1644511149
transform 1 0 94668 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1029
timestamp 1644511149
transform 1 0 95772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1035
timestamp 1644511149
transform 1 0 96324 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1037
timestamp 1644511149
transform 1 0 96508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1049
timestamp 1644511149
transform 1 0 97612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1061
timestamp 1644511149
transform 1 0 98716 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1073
timestamp 1644511149
transform 1 0 99820 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1085
timestamp 1644511149
transform 1 0 100924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1091
timestamp 1644511149
transform 1 0 101476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1093
timestamp 1644511149
transform 1 0 101660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1105
timestamp 1644511149
transform 1 0 102764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1117
timestamp 1644511149
transform 1 0 103868 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1129
timestamp 1644511149
transform 1 0 104972 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1141
timestamp 1644511149
transform 1 0 106076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1147
timestamp 1644511149
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1149
timestamp 1644511149
transform 1 0 106812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1161
timestamp 1644511149
transform 1 0 107916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1173
timestamp 1644511149
transform 1 0 109020 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1185
timestamp 1644511149
transform 1 0 110124 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1197
timestamp 1644511149
transform 1 0 111228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1203
timestamp 1644511149
transform 1 0 111780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1205
timestamp 1644511149
transform 1 0 111964 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1217
timestamp 1644511149
transform 1 0 113068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1229
timestamp 1644511149
transform 1 0 114172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1241
timestamp 1644511149
transform 1 0 115276 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1253
timestamp 1644511149
transform 1 0 116380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1259
timestamp 1644511149
transform 1 0 116932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1261
timestamp 1644511149
transform 1 0 117116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_1273
timestamp 1644511149
transform 1 0 118220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_741
timestamp 1644511149
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_753
timestamp 1644511149
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_765
timestamp 1644511149
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1644511149
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1644511149
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_785
timestamp 1644511149
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_797
timestamp 1644511149
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_809
timestamp 1644511149
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_821
timestamp 1644511149
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_833
timestamp 1644511149
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_839
timestamp 1644511149
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_841
timestamp 1644511149
transform 1 0 78476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_853
timestamp 1644511149
transform 1 0 79580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_865
timestamp 1644511149
transform 1 0 80684 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_877
timestamp 1644511149
transform 1 0 81788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_889
timestamp 1644511149
transform 1 0 82892 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_895
timestamp 1644511149
transform 1 0 83444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_897
timestamp 1644511149
transform 1 0 83628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_909
timestamp 1644511149
transform 1 0 84732 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_921
timestamp 1644511149
transform 1 0 85836 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_933
timestamp 1644511149
transform 1 0 86940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_945
timestamp 1644511149
transform 1 0 88044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_951
timestamp 1644511149
transform 1 0 88596 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_953
timestamp 1644511149
transform 1 0 88780 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_965
timestamp 1644511149
transform 1 0 89884 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_977
timestamp 1644511149
transform 1 0 90988 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_989
timestamp 1644511149
transform 1 0 92092 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1001
timestamp 1644511149
transform 1 0 93196 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1007
timestamp 1644511149
transform 1 0 93748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1009
timestamp 1644511149
transform 1 0 93932 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1021
timestamp 1644511149
transform 1 0 95036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1033
timestamp 1644511149
transform 1 0 96140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1045
timestamp 1644511149
transform 1 0 97244 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1057
timestamp 1644511149
transform 1 0 98348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1063
timestamp 1644511149
transform 1 0 98900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1065
timestamp 1644511149
transform 1 0 99084 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1077
timestamp 1644511149
transform 1 0 100188 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1089
timestamp 1644511149
transform 1 0 101292 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1101
timestamp 1644511149
transform 1 0 102396 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1113
timestamp 1644511149
transform 1 0 103500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1119
timestamp 1644511149
transform 1 0 104052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1121
timestamp 1644511149
transform 1 0 104236 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1133
timestamp 1644511149
transform 1 0 105340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1145
timestamp 1644511149
transform 1 0 106444 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1157
timestamp 1644511149
transform 1 0 107548 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1169
timestamp 1644511149
transform 1 0 108652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1175
timestamp 1644511149
transform 1 0 109204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1177
timestamp 1644511149
transform 1 0 109388 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1189
timestamp 1644511149
transform 1 0 110492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1201
timestamp 1644511149
transform 1 0 111596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1213
timestamp 1644511149
transform 1 0 112700 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1225
timestamp 1644511149
transform 1 0 113804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1231
timestamp 1644511149
transform 1 0 114356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1233
timestamp 1644511149
transform 1 0 114540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1245
timestamp 1644511149
transform 1 0 115644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1257
timestamp 1644511149
transform 1 0 116748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1269
timestamp 1644511149
transform 1 0 117852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1644511149
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1644511149
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_645
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1644511149
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1644511149
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1644511149
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1644511149
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1644511149
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_737
timestamp 1644511149
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1644511149
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1644511149
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_757
timestamp 1644511149
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_769
timestamp 1644511149
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_781
timestamp 1644511149
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_793
timestamp 1644511149
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1644511149
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1644511149
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_813
timestamp 1644511149
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_825
timestamp 1644511149
transform 1 0 77004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_837
timestamp 1644511149
transform 1 0 78108 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_849
timestamp 1644511149
transform 1 0 79212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_861
timestamp 1644511149
transform 1 0 80316 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_867
timestamp 1644511149
transform 1 0 80868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_869
timestamp 1644511149
transform 1 0 81052 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_881
timestamp 1644511149
transform 1 0 82156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_893
timestamp 1644511149
transform 1 0 83260 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_905
timestamp 1644511149
transform 1 0 84364 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_917
timestamp 1644511149
transform 1 0 85468 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_923
timestamp 1644511149
transform 1 0 86020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_925
timestamp 1644511149
transform 1 0 86204 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_937
timestamp 1644511149
transform 1 0 87308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_949
timestamp 1644511149
transform 1 0 88412 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_961
timestamp 1644511149
transform 1 0 89516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_973
timestamp 1644511149
transform 1 0 90620 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_979
timestamp 1644511149
transform 1 0 91172 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_981
timestamp 1644511149
transform 1 0 91356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_993
timestamp 1644511149
transform 1 0 92460 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1005
timestamp 1644511149
transform 1 0 93564 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1017
timestamp 1644511149
transform 1 0 94668 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1029
timestamp 1644511149
transform 1 0 95772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1035
timestamp 1644511149
transform 1 0 96324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1037
timestamp 1644511149
transform 1 0 96508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1049
timestamp 1644511149
transform 1 0 97612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1061
timestamp 1644511149
transform 1 0 98716 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1073
timestamp 1644511149
transform 1 0 99820 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1085
timestamp 1644511149
transform 1 0 100924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1091
timestamp 1644511149
transform 1 0 101476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1093
timestamp 1644511149
transform 1 0 101660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1105
timestamp 1644511149
transform 1 0 102764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1117
timestamp 1644511149
transform 1 0 103868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1129
timestamp 1644511149
transform 1 0 104972 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1141
timestamp 1644511149
transform 1 0 106076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1147
timestamp 1644511149
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1149
timestamp 1644511149
transform 1 0 106812 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1161
timestamp 1644511149
transform 1 0 107916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1173
timestamp 1644511149
transform 1 0 109020 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1185
timestamp 1644511149
transform 1 0 110124 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1197
timestamp 1644511149
transform 1 0 111228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1203
timestamp 1644511149
transform 1 0 111780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1205
timestamp 1644511149
transform 1 0 111964 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1217
timestamp 1644511149
transform 1 0 113068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1229
timestamp 1644511149
transform 1 0 114172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1241
timestamp 1644511149
transform 1 0 115276 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1253
timestamp 1644511149
transform 1 0 116380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1259
timestamp 1644511149
transform 1 0 116932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1261
timestamp 1644511149
transform 1 0 117116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1273
timestamp 1644511149
transform 1 0 118220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_629
timestamp 1644511149
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_641
timestamp 1644511149
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_653
timestamp 1644511149
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1644511149
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_741
timestamp 1644511149
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_753
timestamp 1644511149
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_765
timestamp 1644511149
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1644511149
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1644511149
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_785
timestamp 1644511149
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_797
timestamp 1644511149
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_809
timestamp 1644511149
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_821
timestamp 1644511149
transform 1 0 76636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_833
timestamp 1644511149
transform 1 0 77740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_839
timestamp 1644511149
transform 1 0 78292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_841
timestamp 1644511149
transform 1 0 78476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_853
timestamp 1644511149
transform 1 0 79580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_865
timestamp 1644511149
transform 1 0 80684 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_877
timestamp 1644511149
transform 1 0 81788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_889
timestamp 1644511149
transform 1 0 82892 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_895
timestamp 1644511149
transform 1 0 83444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_897
timestamp 1644511149
transform 1 0 83628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_909
timestamp 1644511149
transform 1 0 84732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_921
timestamp 1644511149
transform 1 0 85836 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_933
timestamp 1644511149
transform 1 0 86940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_945
timestamp 1644511149
transform 1 0 88044 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_951
timestamp 1644511149
transform 1 0 88596 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_953
timestamp 1644511149
transform 1 0 88780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_965
timestamp 1644511149
transform 1 0 89884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_977
timestamp 1644511149
transform 1 0 90988 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_989
timestamp 1644511149
transform 1 0 92092 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1001
timestamp 1644511149
transform 1 0 93196 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1007
timestamp 1644511149
transform 1 0 93748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1009
timestamp 1644511149
transform 1 0 93932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1021
timestamp 1644511149
transform 1 0 95036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1033
timestamp 1644511149
transform 1 0 96140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1045
timestamp 1644511149
transform 1 0 97244 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1057
timestamp 1644511149
transform 1 0 98348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1063
timestamp 1644511149
transform 1 0 98900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1065
timestamp 1644511149
transform 1 0 99084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1077
timestamp 1644511149
transform 1 0 100188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1089
timestamp 1644511149
transform 1 0 101292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1101
timestamp 1644511149
transform 1 0 102396 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1113
timestamp 1644511149
transform 1 0 103500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1119
timestamp 1644511149
transform 1 0 104052 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1121
timestamp 1644511149
transform 1 0 104236 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1133
timestamp 1644511149
transform 1 0 105340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1145
timestamp 1644511149
transform 1 0 106444 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1157
timestamp 1644511149
transform 1 0 107548 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1169
timestamp 1644511149
transform 1 0 108652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1175
timestamp 1644511149
transform 1 0 109204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1177
timestamp 1644511149
transform 1 0 109388 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1189
timestamp 1644511149
transform 1 0 110492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1201
timestamp 1644511149
transform 1 0 111596 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1213
timestamp 1644511149
transform 1 0 112700 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1225
timestamp 1644511149
transform 1 0 113804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1231
timestamp 1644511149
transform 1 0 114356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1233
timestamp 1644511149
transform 1 0 114540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1245
timestamp 1644511149
transform 1 0 115644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1257
timestamp 1644511149
transform 1 0 116748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_1269
timestamp 1644511149
transform 1 0 117852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1644511149
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_645
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1644511149
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1644511149
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1644511149
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1644511149
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1644511149
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_737
timestamp 1644511149
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1644511149
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1644511149
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_757
timestamp 1644511149
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_769
timestamp 1644511149
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_781
timestamp 1644511149
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_793
timestamp 1644511149
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1644511149
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1644511149
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_813
timestamp 1644511149
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1644511149
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_837
timestamp 1644511149
transform 1 0 78108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_849
timestamp 1644511149
transform 1 0 79212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_861
timestamp 1644511149
transform 1 0 80316 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_867
timestamp 1644511149
transform 1 0 80868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_869
timestamp 1644511149
transform 1 0 81052 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_881
timestamp 1644511149
transform 1 0 82156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_893
timestamp 1644511149
transform 1 0 83260 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_905
timestamp 1644511149
transform 1 0 84364 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_917
timestamp 1644511149
transform 1 0 85468 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_923
timestamp 1644511149
transform 1 0 86020 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_925
timestamp 1644511149
transform 1 0 86204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_937
timestamp 1644511149
transform 1 0 87308 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_949
timestamp 1644511149
transform 1 0 88412 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_961
timestamp 1644511149
transform 1 0 89516 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_973
timestamp 1644511149
transform 1 0 90620 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_979
timestamp 1644511149
transform 1 0 91172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_981
timestamp 1644511149
transform 1 0 91356 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_993
timestamp 1644511149
transform 1 0 92460 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1005
timestamp 1644511149
transform 1 0 93564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1017
timestamp 1644511149
transform 1 0 94668 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1029
timestamp 1644511149
transform 1 0 95772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1035
timestamp 1644511149
transform 1 0 96324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1037
timestamp 1644511149
transform 1 0 96508 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1049
timestamp 1644511149
transform 1 0 97612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1061
timestamp 1644511149
transform 1 0 98716 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1073
timestamp 1644511149
transform 1 0 99820 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1085
timestamp 1644511149
transform 1 0 100924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1091
timestamp 1644511149
transform 1 0 101476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1093
timestamp 1644511149
transform 1 0 101660 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1105
timestamp 1644511149
transform 1 0 102764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1117
timestamp 1644511149
transform 1 0 103868 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1129
timestamp 1644511149
transform 1 0 104972 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1141
timestamp 1644511149
transform 1 0 106076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1147
timestamp 1644511149
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1149
timestamp 1644511149
transform 1 0 106812 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1161
timestamp 1644511149
transform 1 0 107916 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1173
timestamp 1644511149
transform 1 0 109020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1185
timestamp 1644511149
transform 1 0 110124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1197
timestamp 1644511149
transform 1 0 111228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1203
timestamp 1644511149
transform 1 0 111780 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1205
timestamp 1644511149
transform 1 0 111964 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1217
timestamp 1644511149
transform 1 0 113068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1229
timestamp 1644511149
transform 1 0 114172 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1241
timestamp 1644511149
transform 1 0 115276 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1253
timestamp 1644511149
transform 1 0 116380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1259
timestamp 1644511149
transform 1 0 116932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1261
timestamp 1644511149
transform 1 0 117116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_1273
timestamp 1644511149
transform 1 0 118220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1644511149
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1644511149
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1644511149
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1644511149
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1644511149
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1644511149
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1644511149
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_741
timestamp 1644511149
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_753
timestamp 1644511149
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_765
timestamp 1644511149
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1644511149
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1644511149
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_785
timestamp 1644511149
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_797
timestamp 1644511149
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_809
timestamp 1644511149
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_821
timestamp 1644511149
transform 1 0 76636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_833
timestamp 1644511149
transform 1 0 77740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_839
timestamp 1644511149
transform 1 0 78292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_841
timestamp 1644511149
transform 1 0 78476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_853
timestamp 1644511149
transform 1 0 79580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_865
timestamp 1644511149
transform 1 0 80684 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_877
timestamp 1644511149
transform 1 0 81788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_889
timestamp 1644511149
transform 1 0 82892 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_895
timestamp 1644511149
transform 1 0 83444 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_897
timestamp 1644511149
transform 1 0 83628 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_909
timestamp 1644511149
transform 1 0 84732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_921
timestamp 1644511149
transform 1 0 85836 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_933
timestamp 1644511149
transform 1 0 86940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_945
timestamp 1644511149
transform 1 0 88044 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_951
timestamp 1644511149
transform 1 0 88596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_953
timestamp 1644511149
transform 1 0 88780 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_965
timestamp 1644511149
transform 1 0 89884 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_977
timestamp 1644511149
transform 1 0 90988 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_989
timestamp 1644511149
transform 1 0 92092 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1001
timestamp 1644511149
transform 1 0 93196 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1007
timestamp 1644511149
transform 1 0 93748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1009
timestamp 1644511149
transform 1 0 93932 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1021
timestamp 1644511149
transform 1 0 95036 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1033
timestamp 1644511149
transform 1 0 96140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1045
timestamp 1644511149
transform 1 0 97244 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1057
timestamp 1644511149
transform 1 0 98348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1063
timestamp 1644511149
transform 1 0 98900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1065
timestamp 1644511149
transform 1 0 99084 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1077
timestamp 1644511149
transform 1 0 100188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1089
timestamp 1644511149
transform 1 0 101292 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1101
timestamp 1644511149
transform 1 0 102396 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1113
timestamp 1644511149
transform 1 0 103500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1119
timestamp 1644511149
transform 1 0 104052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1121
timestamp 1644511149
transform 1 0 104236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1133
timestamp 1644511149
transform 1 0 105340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1145
timestamp 1644511149
transform 1 0 106444 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1157
timestamp 1644511149
transform 1 0 107548 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1169
timestamp 1644511149
transform 1 0 108652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1175
timestamp 1644511149
transform 1 0 109204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1177
timestamp 1644511149
transform 1 0 109388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1189
timestamp 1644511149
transform 1 0 110492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1201
timestamp 1644511149
transform 1 0 111596 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1213
timestamp 1644511149
transform 1 0 112700 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1225
timestamp 1644511149
transform 1 0 113804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1231
timestamp 1644511149
transform 1 0 114356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1233
timestamp 1644511149
transform 1 0 114540 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1245
timestamp 1644511149
transform 1 0 115644 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1257
timestamp 1644511149
transform 1 0 116748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_1269
timestamp 1644511149
transform 1 0 117852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1644511149
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1644511149
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1644511149
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_701
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_713
timestamp 1644511149
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_725
timestamp 1644511149
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_737
timestamp 1644511149
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1644511149
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1644511149
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_757
timestamp 1644511149
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_769
timestamp 1644511149
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_781
timestamp 1644511149
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_793
timestamp 1644511149
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1644511149
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1644511149
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_813
timestamp 1644511149
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_825
timestamp 1644511149
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_837
timestamp 1644511149
transform 1 0 78108 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_849
timestamp 1644511149
transform 1 0 79212 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_861
timestamp 1644511149
transform 1 0 80316 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_867
timestamp 1644511149
transform 1 0 80868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_869
timestamp 1644511149
transform 1 0 81052 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_881
timestamp 1644511149
transform 1 0 82156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_893
timestamp 1644511149
transform 1 0 83260 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_905
timestamp 1644511149
transform 1 0 84364 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_917
timestamp 1644511149
transform 1 0 85468 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_923
timestamp 1644511149
transform 1 0 86020 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_925
timestamp 1644511149
transform 1 0 86204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_937
timestamp 1644511149
transform 1 0 87308 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_949
timestamp 1644511149
transform 1 0 88412 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_961
timestamp 1644511149
transform 1 0 89516 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_973
timestamp 1644511149
transform 1 0 90620 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_979
timestamp 1644511149
transform 1 0 91172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_981
timestamp 1644511149
transform 1 0 91356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_993
timestamp 1644511149
transform 1 0 92460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1005
timestamp 1644511149
transform 1 0 93564 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1017
timestamp 1644511149
transform 1 0 94668 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1029
timestamp 1644511149
transform 1 0 95772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1035
timestamp 1644511149
transform 1 0 96324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1037
timestamp 1644511149
transform 1 0 96508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1049
timestamp 1644511149
transform 1 0 97612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1061
timestamp 1644511149
transform 1 0 98716 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1073
timestamp 1644511149
transform 1 0 99820 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1085
timestamp 1644511149
transform 1 0 100924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1091
timestamp 1644511149
transform 1 0 101476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1093
timestamp 1644511149
transform 1 0 101660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1105
timestamp 1644511149
transform 1 0 102764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1117
timestamp 1644511149
transform 1 0 103868 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1129
timestamp 1644511149
transform 1 0 104972 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1141
timestamp 1644511149
transform 1 0 106076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1147
timestamp 1644511149
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1149
timestamp 1644511149
transform 1 0 106812 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1161
timestamp 1644511149
transform 1 0 107916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1173
timestamp 1644511149
transform 1 0 109020 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1185
timestamp 1644511149
transform 1 0 110124 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1197
timestamp 1644511149
transform 1 0 111228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1203
timestamp 1644511149
transform 1 0 111780 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1205
timestamp 1644511149
transform 1 0 111964 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1217
timestamp 1644511149
transform 1 0 113068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1229
timestamp 1644511149
transform 1 0 114172 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1241
timestamp 1644511149
transform 1 0 115276 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1253
timestamp 1644511149
transform 1 0 116380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1259
timestamp 1644511149
transform 1 0 116932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1261
timestamp 1644511149
transform 1 0 117116 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1273
timestamp 1644511149
transform 1 0 118220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1644511149
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1644511149
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1644511149
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_741
timestamp 1644511149
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_753
timestamp 1644511149
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_765
timestamp 1644511149
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1644511149
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1644511149
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_785
timestamp 1644511149
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_797
timestamp 1644511149
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_809
timestamp 1644511149
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_821
timestamp 1644511149
transform 1 0 76636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_833
timestamp 1644511149
transform 1 0 77740 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_839
timestamp 1644511149
transform 1 0 78292 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_841
timestamp 1644511149
transform 1 0 78476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_853
timestamp 1644511149
transform 1 0 79580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_865
timestamp 1644511149
transform 1 0 80684 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_877
timestamp 1644511149
transform 1 0 81788 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_889
timestamp 1644511149
transform 1 0 82892 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_895
timestamp 1644511149
transform 1 0 83444 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_897
timestamp 1644511149
transform 1 0 83628 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_909
timestamp 1644511149
transform 1 0 84732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_921
timestamp 1644511149
transform 1 0 85836 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_933
timestamp 1644511149
transform 1 0 86940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_945
timestamp 1644511149
transform 1 0 88044 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_951
timestamp 1644511149
transform 1 0 88596 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_953
timestamp 1644511149
transform 1 0 88780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_965
timestamp 1644511149
transform 1 0 89884 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_977
timestamp 1644511149
transform 1 0 90988 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_989
timestamp 1644511149
transform 1 0 92092 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1001
timestamp 1644511149
transform 1 0 93196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1007
timestamp 1644511149
transform 1 0 93748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1009
timestamp 1644511149
transform 1 0 93932 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1021
timestamp 1644511149
transform 1 0 95036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1033
timestamp 1644511149
transform 1 0 96140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1045
timestamp 1644511149
transform 1 0 97244 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1057
timestamp 1644511149
transform 1 0 98348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1063
timestamp 1644511149
transform 1 0 98900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1065
timestamp 1644511149
transform 1 0 99084 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1077
timestamp 1644511149
transform 1 0 100188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1089
timestamp 1644511149
transform 1 0 101292 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1101
timestamp 1644511149
transform 1 0 102396 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1113
timestamp 1644511149
transform 1 0 103500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1119
timestamp 1644511149
transform 1 0 104052 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1121
timestamp 1644511149
transform 1 0 104236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1133
timestamp 1644511149
transform 1 0 105340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1145
timestamp 1644511149
transform 1 0 106444 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1157
timestamp 1644511149
transform 1 0 107548 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1169
timestamp 1644511149
transform 1 0 108652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1175
timestamp 1644511149
transform 1 0 109204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1177
timestamp 1644511149
transform 1 0 109388 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1189
timestamp 1644511149
transform 1 0 110492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1201
timestamp 1644511149
transform 1 0 111596 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1213
timestamp 1644511149
transform 1 0 112700 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1225
timestamp 1644511149
transform 1 0 113804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1231
timestamp 1644511149
transform 1 0 114356 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1233
timestamp 1644511149
transform 1 0 114540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1245
timestamp 1644511149
transform 1 0 115644 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1257
timestamp 1644511149
transform 1 0 116748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_1269
timestamp 1644511149
transform 1 0 117852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_625
timestamp 1644511149
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1644511149
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1644511149
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_713
timestamp 1644511149
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_725
timestamp 1644511149
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_737
timestamp 1644511149
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1644511149
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1644511149
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_757
timestamp 1644511149
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_769
timestamp 1644511149
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_781
timestamp 1644511149
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_793
timestamp 1644511149
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1644511149
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1644511149
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_813
timestamp 1644511149
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_825
timestamp 1644511149
transform 1 0 77004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_837
timestamp 1644511149
transform 1 0 78108 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_849
timestamp 1644511149
transform 1 0 79212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_861
timestamp 1644511149
transform 1 0 80316 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_867
timestamp 1644511149
transform 1 0 80868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_869
timestamp 1644511149
transform 1 0 81052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_881
timestamp 1644511149
transform 1 0 82156 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_893
timestamp 1644511149
transform 1 0 83260 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_905
timestamp 1644511149
transform 1 0 84364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_917
timestamp 1644511149
transform 1 0 85468 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_923
timestamp 1644511149
transform 1 0 86020 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_925
timestamp 1644511149
transform 1 0 86204 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_937
timestamp 1644511149
transform 1 0 87308 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_949
timestamp 1644511149
transform 1 0 88412 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_961
timestamp 1644511149
transform 1 0 89516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_973
timestamp 1644511149
transform 1 0 90620 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_979
timestamp 1644511149
transform 1 0 91172 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_981
timestamp 1644511149
transform 1 0 91356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_993
timestamp 1644511149
transform 1 0 92460 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1005
timestamp 1644511149
transform 1 0 93564 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1017
timestamp 1644511149
transform 1 0 94668 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1029
timestamp 1644511149
transform 1 0 95772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1035
timestamp 1644511149
transform 1 0 96324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1037
timestamp 1644511149
transform 1 0 96508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1049
timestamp 1644511149
transform 1 0 97612 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1061
timestamp 1644511149
transform 1 0 98716 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1073
timestamp 1644511149
transform 1 0 99820 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1085
timestamp 1644511149
transform 1 0 100924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1091
timestamp 1644511149
transform 1 0 101476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1093
timestamp 1644511149
transform 1 0 101660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1105
timestamp 1644511149
transform 1 0 102764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1117
timestamp 1644511149
transform 1 0 103868 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1129
timestamp 1644511149
transform 1 0 104972 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1141
timestamp 1644511149
transform 1 0 106076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1147
timestamp 1644511149
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1149
timestamp 1644511149
transform 1 0 106812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1161
timestamp 1644511149
transform 1 0 107916 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1173
timestamp 1644511149
transform 1 0 109020 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1185
timestamp 1644511149
transform 1 0 110124 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1197
timestamp 1644511149
transform 1 0 111228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1203
timestamp 1644511149
transform 1 0 111780 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1205
timestamp 1644511149
transform 1 0 111964 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1217
timestamp 1644511149
transform 1 0 113068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1229
timestamp 1644511149
transform 1 0 114172 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1241
timestamp 1644511149
transform 1 0 115276 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1253
timestamp 1644511149
transform 1 0 116380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1259
timestamp 1644511149
transform 1 0 116932 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1261
timestamp 1644511149
transform 1 0 117116 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_1273
timestamp 1644511149
transform 1 0 118220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1644511149
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_741
timestamp 1644511149
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_753
timestamp 1644511149
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_765
timestamp 1644511149
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1644511149
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1644511149
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_785
timestamp 1644511149
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_797
timestamp 1644511149
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_809
timestamp 1644511149
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_821
timestamp 1644511149
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_833
timestamp 1644511149
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_839
timestamp 1644511149
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_841
timestamp 1644511149
transform 1 0 78476 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_853
timestamp 1644511149
transform 1 0 79580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_865
timestamp 1644511149
transform 1 0 80684 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_877
timestamp 1644511149
transform 1 0 81788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_889
timestamp 1644511149
transform 1 0 82892 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_895
timestamp 1644511149
transform 1 0 83444 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_897
timestamp 1644511149
transform 1 0 83628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_909
timestamp 1644511149
transform 1 0 84732 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_921
timestamp 1644511149
transform 1 0 85836 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_933
timestamp 1644511149
transform 1 0 86940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_945
timestamp 1644511149
transform 1 0 88044 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_951
timestamp 1644511149
transform 1 0 88596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_953
timestamp 1644511149
transform 1 0 88780 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_965
timestamp 1644511149
transform 1 0 89884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_977
timestamp 1644511149
transform 1 0 90988 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_989
timestamp 1644511149
transform 1 0 92092 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1001
timestamp 1644511149
transform 1 0 93196 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1007
timestamp 1644511149
transform 1 0 93748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1009
timestamp 1644511149
transform 1 0 93932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1021
timestamp 1644511149
transform 1 0 95036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1033
timestamp 1644511149
transform 1 0 96140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1045
timestamp 1644511149
transform 1 0 97244 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1057
timestamp 1644511149
transform 1 0 98348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1063
timestamp 1644511149
transform 1 0 98900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1065
timestamp 1644511149
transform 1 0 99084 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1077
timestamp 1644511149
transform 1 0 100188 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1089
timestamp 1644511149
transform 1 0 101292 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1101
timestamp 1644511149
transform 1 0 102396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1113
timestamp 1644511149
transform 1 0 103500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1119
timestamp 1644511149
transform 1 0 104052 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1121
timestamp 1644511149
transform 1 0 104236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1133
timestamp 1644511149
transform 1 0 105340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1145
timestamp 1644511149
transform 1 0 106444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1157
timestamp 1644511149
transform 1 0 107548 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1169
timestamp 1644511149
transform 1 0 108652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1175
timestamp 1644511149
transform 1 0 109204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1177
timestamp 1644511149
transform 1 0 109388 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1189
timestamp 1644511149
transform 1 0 110492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1201
timestamp 1644511149
transform 1 0 111596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1213
timestamp 1644511149
transform 1 0 112700 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1225
timestamp 1644511149
transform 1 0 113804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1231
timestamp 1644511149
transform 1 0 114356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1233
timestamp 1644511149
transform 1 0 114540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1245
timestamp 1644511149
transform 1 0 115644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1257
timestamp 1644511149
transform 1 0 116748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_1269
timestamp 1644511149
transform 1 0 117852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_625
timestamp 1644511149
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1644511149
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1644511149
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_725
timestamp 1644511149
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_737
timestamp 1644511149
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 1644511149
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1644511149
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_757
timestamp 1644511149
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_769
timestamp 1644511149
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_781
timestamp 1644511149
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_793
timestamp 1644511149
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1644511149
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1644511149
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_813
timestamp 1644511149
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_825
timestamp 1644511149
transform 1 0 77004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_837
timestamp 1644511149
transform 1 0 78108 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_849
timestamp 1644511149
transform 1 0 79212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_861
timestamp 1644511149
transform 1 0 80316 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_867
timestamp 1644511149
transform 1 0 80868 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_869
timestamp 1644511149
transform 1 0 81052 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_881
timestamp 1644511149
transform 1 0 82156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_893
timestamp 1644511149
transform 1 0 83260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_905
timestamp 1644511149
transform 1 0 84364 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_917
timestamp 1644511149
transform 1 0 85468 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_923
timestamp 1644511149
transform 1 0 86020 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_925
timestamp 1644511149
transform 1 0 86204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_937
timestamp 1644511149
transform 1 0 87308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_949
timestamp 1644511149
transform 1 0 88412 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_961
timestamp 1644511149
transform 1 0 89516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_973
timestamp 1644511149
transform 1 0 90620 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_979
timestamp 1644511149
transform 1 0 91172 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_981
timestamp 1644511149
transform 1 0 91356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_993
timestamp 1644511149
transform 1 0 92460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1005
timestamp 1644511149
transform 1 0 93564 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1017
timestamp 1644511149
transform 1 0 94668 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1029
timestamp 1644511149
transform 1 0 95772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1035
timestamp 1644511149
transform 1 0 96324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1037
timestamp 1644511149
transform 1 0 96508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1049
timestamp 1644511149
transform 1 0 97612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1061
timestamp 1644511149
transform 1 0 98716 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1073
timestamp 1644511149
transform 1 0 99820 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1085
timestamp 1644511149
transform 1 0 100924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1091
timestamp 1644511149
transform 1 0 101476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1093
timestamp 1644511149
transform 1 0 101660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1105
timestamp 1644511149
transform 1 0 102764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1117
timestamp 1644511149
transform 1 0 103868 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1129
timestamp 1644511149
transform 1 0 104972 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1141
timestamp 1644511149
transform 1 0 106076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1147
timestamp 1644511149
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1149
timestamp 1644511149
transform 1 0 106812 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1161
timestamp 1644511149
transform 1 0 107916 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1173
timestamp 1644511149
transform 1 0 109020 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1185
timestamp 1644511149
transform 1 0 110124 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1197
timestamp 1644511149
transform 1 0 111228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1203
timestamp 1644511149
transform 1 0 111780 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1205
timestamp 1644511149
transform 1 0 111964 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1217
timestamp 1644511149
transform 1 0 113068 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1229
timestamp 1644511149
transform 1 0 114172 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1241
timestamp 1644511149
transform 1 0 115276 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1253
timestamp 1644511149
transform 1 0 116380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1259
timestamp 1644511149
transform 1 0 116932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1261
timestamp 1644511149
transform 1 0 117116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_1267
timestamp 1644511149
transform 1 0 117668 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1273
timestamp 1644511149
transform 1 0 118220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_19
timestamp 1644511149
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_31
timestamp 1644511149
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_43
timestamp 1644511149
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1644511149
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1644511149
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_741
timestamp 1644511149
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_753
timestamp 1644511149
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_765
timestamp 1644511149
transform 1 0 71484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 1644511149
transform 1 0 72588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 1644511149
transform 1 0 73140 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_785
timestamp 1644511149
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_797
timestamp 1644511149
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_809
timestamp 1644511149
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_821
timestamp 1644511149
transform 1 0 76636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_833
timestamp 1644511149
transform 1 0 77740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_839
timestamp 1644511149
transform 1 0 78292 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_841
timestamp 1644511149
transform 1 0 78476 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_853
timestamp 1644511149
transform 1 0 79580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_865
timestamp 1644511149
transform 1 0 80684 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_877
timestamp 1644511149
transform 1 0 81788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_889
timestamp 1644511149
transform 1 0 82892 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_895
timestamp 1644511149
transform 1 0 83444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_897
timestamp 1644511149
transform 1 0 83628 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_909
timestamp 1644511149
transform 1 0 84732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_921
timestamp 1644511149
transform 1 0 85836 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_933
timestamp 1644511149
transform 1 0 86940 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_945
timestamp 1644511149
transform 1 0 88044 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_951
timestamp 1644511149
transform 1 0 88596 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_953
timestamp 1644511149
transform 1 0 88780 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_965
timestamp 1644511149
transform 1 0 89884 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_977
timestamp 1644511149
transform 1 0 90988 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_989
timestamp 1644511149
transform 1 0 92092 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1001
timestamp 1644511149
transform 1 0 93196 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1007
timestamp 1644511149
transform 1 0 93748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1009
timestamp 1644511149
transform 1 0 93932 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1021
timestamp 1644511149
transform 1 0 95036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1033
timestamp 1644511149
transform 1 0 96140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1045
timestamp 1644511149
transform 1 0 97244 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1057
timestamp 1644511149
transform 1 0 98348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1063
timestamp 1644511149
transform 1 0 98900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1065
timestamp 1644511149
transform 1 0 99084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1077
timestamp 1644511149
transform 1 0 100188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1089
timestamp 1644511149
transform 1 0 101292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1101
timestamp 1644511149
transform 1 0 102396 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1113
timestamp 1644511149
transform 1 0 103500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1119
timestamp 1644511149
transform 1 0 104052 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1121
timestamp 1644511149
transform 1 0 104236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1133
timestamp 1644511149
transform 1 0 105340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1145
timestamp 1644511149
transform 1 0 106444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1157
timestamp 1644511149
transform 1 0 107548 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1169
timestamp 1644511149
transform 1 0 108652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1175
timestamp 1644511149
transform 1 0 109204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1177
timestamp 1644511149
transform 1 0 109388 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1189
timestamp 1644511149
transform 1 0 110492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1201
timestamp 1644511149
transform 1 0 111596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1213
timestamp 1644511149
transform 1 0 112700 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1225
timestamp 1644511149
transform 1 0 113804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1231
timestamp 1644511149
transform 1 0 114356 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1233
timestamp 1644511149
transform 1 0 114540 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1245
timestamp 1644511149
transform 1 0 115644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1257
timestamp 1644511149
transform 1 0 116748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1269
timestamp 1644511149
transform 1 0 117852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_725
timestamp 1644511149
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_737
timestamp 1644511149
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 1644511149
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 1644511149
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_757
timestamp 1644511149
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_769
timestamp 1644511149
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_781
timestamp 1644511149
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_793
timestamp 1644511149
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1644511149
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1644511149
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_813
timestamp 1644511149
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_825
timestamp 1644511149
transform 1 0 77004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_837
timestamp 1644511149
transform 1 0 78108 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_849
timestamp 1644511149
transform 1 0 79212 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_861
timestamp 1644511149
transform 1 0 80316 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_867
timestamp 1644511149
transform 1 0 80868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_869
timestamp 1644511149
transform 1 0 81052 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_881
timestamp 1644511149
transform 1 0 82156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_893
timestamp 1644511149
transform 1 0 83260 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_905
timestamp 1644511149
transform 1 0 84364 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_917
timestamp 1644511149
transform 1 0 85468 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_923
timestamp 1644511149
transform 1 0 86020 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_925
timestamp 1644511149
transform 1 0 86204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_937
timestamp 1644511149
transform 1 0 87308 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_949
timestamp 1644511149
transform 1 0 88412 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_961
timestamp 1644511149
transform 1 0 89516 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_973
timestamp 1644511149
transform 1 0 90620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_979
timestamp 1644511149
transform 1 0 91172 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_981
timestamp 1644511149
transform 1 0 91356 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_993
timestamp 1644511149
transform 1 0 92460 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1005
timestamp 1644511149
transform 1 0 93564 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1017
timestamp 1644511149
transform 1 0 94668 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1029
timestamp 1644511149
transform 1 0 95772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1035
timestamp 1644511149
transform 1 0 96324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1037
timestamp 1644511149
transform 1 0 96508 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1049
timestamp 1644511149
transform 1 0 97612 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1061
timestamp 1644511149
transform 1 0 98716 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1073
timestamp 1644511149
transform 1 0 99820 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1085
timestamp 1644511149
transform 1 0 100924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1091
timestamp 1644511149
transform 1 0 101476 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1093
timestamp 1644511149
transform 1 0 101660 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1105
timestamp 1644511149
transform 1 0 102764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1117
timestamp 1644511149
transform 1 0 103868 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1129
timestamp 1644511149
transform 1 0 104972 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1141
timestamp 1644511149
transform 1 0 106076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1147
timestamp 1644511149
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1149
timestamp 1644511149
transform 1 0 106812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1161
timestamp 1644511149
transform 1 0 107916 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1173
timestamp 1644511149
transform 1 0 109020 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1185
timestamp 1644511149
transform 1 0 110124 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1197
timestamp 1644511149
transform 1 0 111228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1203
timestamp 1644511149
transform 1 0 111780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1205
timestamp 1644511149
transform 1 0 111964 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1217
timestamp 1644511149
transform 1 0 113068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1229
timestamp 1644511149
transform 1 0 114172 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1241
timestamp 1644511149
transform 1 0 115276 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1253
timestamp 1644511149
transform 1 0 116380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1259
timestamp 1644511149
transform 1 0 116932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1261
timestamp 1644511149
transform 1 0 117116 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_1267
timestamp 1644511149
transform 1 0 117668 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1273
timestamp 1644511149
transform 1 0 118220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1644511149
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1644511149
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1644511149
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_741
timestamp 1644511149
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_753
timestamp 1644511149
transform 1 0 70380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_765
timestamp 1644511149
transform 1 0 71484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 1644511149
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 1644511149
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_785
timestamp 1644511149
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_797
timestamp 1644511149
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_809
timestamp 1644511149
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_821
timestamp 1644511149
transform 1 0 76636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_833
timestamp 1644511149
transform 1 0 77740 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_839
timestamp 1644511149
transform 1 0 78292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_841
timestamp 1644511149
transform 1 0 78476 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_853
timestamp 1644511149
transform 1 0 79580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_865
timestamp 1644511149
transform 1 0 80684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_877
timestamp 1644511149
transform 1 0 81788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_889
timestamp 1644511149
transform 1 0 82892 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_895
timestamp 1644511149
transform 1 0 83444 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_897
timestamp 1644511149
transform 1 0 83628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_909
timestamp 1644511149
transform 1 0 84732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_921
timestamp 1644511149
transform 1 0 85836 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_933
timestamp 1644511149
transform 1 0 86940 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_945
timestamp 1644511149
transform 1 0 88044 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_951
timestamp 1644511149
transform 1 0 88596 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_953
timestamp 1644511149
transform 1 0 88780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_965
timestamp 1644511149
transform 1 0 89884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_977
timestamp 1644511149
transform 1 0 90988 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_989
timestamp 1644511149
transform 1 0 92092 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1001
timestamp 1644511149
transform 1 0 93196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1007
timestamp 1644511149
transform 1 0 93748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1009
timestamp 1644511149
transform 1 0 93932 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1021
timestamp 1644511149
transform 1 0 95036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1033
timestamp 1644511149
transform 1 0 96140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1045
timestamp 1644511149
transform 1 0 97244 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1057
timestamp 1644511149
transform 1 0 98348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1063
timestamp 1644511149
transform 1 0 98900 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1065
timestamp 1644511149
transform 1 0 99084 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1077
timestamp 1644511149
transform 1 0 100188 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1089
timestamp 1644511149
transform 1 0 101292 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1101
timestamp 1644511149
transform 1 0 102396 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1113
timestamp 1644511149
transform 1 0 103500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1119
timestamp 1644511149
transform 1 0 104052 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1121
timestamp 1644511149
transform 1 0 104236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1133
timestamp 1644511149
transform 1 0 105340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1145
timestamp 1644511149
transform 1 0 106444 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1157
timestamp 1644511149
transform 1 0 107548 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1169
timestamp 1644511149
transform 1 0 108652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1175
timestamp 1644511149
transform 1 0 109204 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1177
timestamp 1644511149
transform 1 0 109388 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1189
timestamp 1644511149
transform 1 0 110492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1201
timestamp 1644511149
transform 1 0 111596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1213
timestamp 1644511149
transform 1 0 112700 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1225
timestamp 1644511149
transform 1 0 113804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1231
timestamp 1644511149
transform 1 0 114356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1233
timestamp 1644511149
transform 1 0 114540 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1245
timestamp 1644511149
transform 1 0 115644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1257
timestamp 1644511149
transform 1 0 116748 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1269
timestamp 1644511149
transform 1 0 117852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_12
timestamp 1644511149
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_713
timestamp 1644511149
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_725
timestamp 1644511149
transform 1 0 67804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_737
timestamp 1644511149
transform 1 0 68908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1644511149
transform 1 0 70012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1644511149
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_757
timestamp 1644511149
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_769
timestamp 1644511149
transform 1 0 71852 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_781
timestamp 1644511149
transform 1 0 72956 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_793
timestamp 1644511149
transform 1 0 74060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 1644511149
transform 1 0 75164 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1644511149
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_813
timestamp 1644511149
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_825
timestamp 1644511149
transform 1 0 77004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_837
timestamp 1644511149
transform 1 0 78108 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_849
timestamp 1644511149
transform 1 0 79212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_861
timestamp 1644511149
transform 1 0 80316 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_867
timestamp 1644511149
transform 1 0 80868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_869
timestamp 1644511149
transform 1 0 81052 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_881
timestamp 1644511149
transform 1 0 82156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_893
timestamp 1644511149
transform 1 0 83260 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_905
timestamp 1644511149
transform 1 0 84364 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_917
timestamp 1644511149
transform 1 0 85468 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_923
timestamp 1644511149
transform 1 0 86020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_925
timestamp 1644511149
transform 1 0 86204 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_937
timestamp 1644511149
transform 1 0 87308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_949
timestamp 1644511149
transform 1 0 88412 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_961
timestamp 1644511149
transform 1 0 89516 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_973
timestamp 1644511149
transform 1 0 90620 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_979
timestamp 1644511149
transform 1 0 91172 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_981
timestamp 1644511149
transform 1 0 91356 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_993
timestamp 1644511149
transform 1 0 92460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1005
timestamp 1644511149
transform 1 0 93564 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1017
timestamp 1644511149
transform 1 0 94668 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1029
timestamp 1644511149
transform 1 0 95772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1035
timestamp 1644511149
transform 1 0 96324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1037
timestamp 1644511149
transform 1 0 96508 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1049
timestamp 1644511149
transform 1 0 97612 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1061
timestamp 1644511149
transform 1 0 98716 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1073
timestamp 1644511149
transform 1 0 99820 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1085
timestamp 1644511149
transform 1 0 100924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1091
timestamp 1644511149
transform 1 0 101476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1093
timestamp 1644511149
transform 1 0 101660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1105
timestamp 1644511149
transform 1 0 102764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1117
timestamp 1644511149
transform 1 0 103868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1129
timestamp 1644511149
transform 1 0 104972 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1141
timestamp 1644511149
transform 1 0 106076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1147
timestamp 1644511149
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1149
timestamp 1644511149
transform 1 0 106812 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1161
timestamp 1644511149
transform 1 0 107916 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1173
timestamp 1644511149
transform 1 0 109020 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1185
timestamp 1644511149
transform 1 0 110124 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1197
timestamp 1644511149
transform 1 0 111228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1203
timestamp 1644511149
transform 1 0 111780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1205
timestamp 1644511149
transform 1 0 111964 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1217
timestamp 1644511149
transform 1 0 113068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1229
timestamp 1644511149
transform 1 0 114172 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1241
timestamp 1644511149
transform 1 0 115276 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1253
timestamp 1644511149
transform 1 0 116380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1259
timestamp 1644511149
transform 1 0 116932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1261
timestamp 1644511149
transform 1 0 117116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1273
timestamp 1644511149
transform 1 0 118220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_11
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_23
timestamp 1644511149
transform 1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1644511149
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1644511149
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1644511149
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1644511149
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_741
timestamp 1644511149
transform 1 0 69276 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_753
timestamp 1644511149
transform 1 0 70380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_765
timestamp 1644511149
transform 1 0 71484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1644511149
transform 1 0 72588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1644511149
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_785
timestamp 1644511149
transform 1 0 73324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_797
timestamp 1644511149
transform 1 0 74428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_809
timestamp 1644511149
transform 1 0 75532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_821
timestamp 1644511149
transform 1 0 76636 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_833
timestamp 1644511149
transform 1 0 77740 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_839
timestamp 1644511149
transform 1 0 78292 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_841
timestamp 1644511149
transform 1 0 78476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_853
timestamp 1644511149
transform 1 0 79580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_865
timestamp 1644511149
transform 1 0 80684 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_877
timestamp 1644511149
transform 1 0 81788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_889
timestamp 1644511149
transform 1 0 82892 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_895
timestamp 1644511149
transform 1 0 83444 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_897
timestamp 1644511149
transform 1 0 83628 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_909
timestamp 1644511149
transform 1 0 84732 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_921
timestamp 1644511149
transform 1 0 85836 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_933
timestamp 1644511149
transform 1 0 86940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_945
timestamp 1644511149
transform 1 0 88044 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_951
timestamp 1644511149
transform 1 0 88596 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_953
timestamp 1644511149
transform 1 0 88780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_965
timestamp 1644511149
transform 1 0 89884 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_977
timestamp 1644511149
transform 1 0 90988 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_989
timestamp 1644511149
transform 1 0 92092 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1001
timestamp 1644511149
transform 1 0 93196 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1007
timestamp 1644511149
transform 1 0 93748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1009
timestamp 1644511149
transform 1 0 93932 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1021
timestamp 1644511149
transform 1 0 95036 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1033
timestamp 1644511149
transform 1 0 96140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1045
timestamp 1644511149
transform 1 0 97244 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1057
timestamp 1644511149
transform 1 0 98348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1063
timestamp 1644511149
transform 1 0 98900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1065
timestamp 1644511149
transform 1 0 99084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1077
timestamp 1644511149
transform 1 0 100188 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1089
timestamp 1644511149
transform 1 0 101292 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1101
timestamp 1644511149
transform 1 0 102396 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1113
timestamp 1644511149
transform 1 0 103500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1119
timestamp 1644511149
transform 1 0 104052 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1121
timestamp 1644511149
transform 1 0 104236 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1133
timestamp 1644511149
transform 1 0 105340 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1145
timestamp 1644511149
transform 1 0 106444 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1157
timestamp 1644511149
transform 1 0 107548 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1169
timestamp 1644511149
transform 1 0 108652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1175
timestamp 1644511149
transform 1 0 109204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1177
timestamp 1644511149
transform 1 0 109388 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1189
timestamp 1644511149
transform 1 0 110492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1201
timestamp 1644511149
transform 1 0 111596 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1213
timestamp 1644511149
transform 1 0 112700 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1225
timestamp 1644511149
transform 1 0 113804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1231
timestamp 1644511149
transform 1 0 114356 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1233
timestamp 1644511149
transform 1 0 114540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1245
timestamp 1644511149
transform 1 0 115644 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1257
timestamp 1644511149
transform 1 0 116748 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1267
timestamp 1644511149
transform 1 0 117668 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1273
timestamp 1644511149
transform 1 0 118220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_19
timestamp 1644511149
transform 1 0 2852 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1644511149
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_103
timestamp 1644511149
transform 1 0 10580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1644511149
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_148
timestamp 1644511149
transform 1 0 14720 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1644511149
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_238
timestamp 1644511149
transform 1 0 23000 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1644511149
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_284
timestamp 1644511149
transform 1 0 27232 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_296
timestamp 1644511149
transform 1 0 28336 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1644511149
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_369
timestamp 1644511149
transform 1 0 35052 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1644511149
transform 1 0 35420 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1644511149
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1644511149
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_405
timestamp 1644511149
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1644511149
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_430
timestamp 1644511149
transform 1 0 40664 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_442
timestamp 1644511149
transform 1 0 41768 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_449
timestamp 1644511149
transform 1 0 42412 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_461
timestamp 1644511149
transform 1 0 43516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_473
timestamp 1644511149
transform 1 0 44620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_509
timestamp 1644511149
transform 1 0 47932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_521
timestamp 1644511149
transform 1 0 49036 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_529
timestamp 1644511149
transform 1 0 49772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_549
timestamp 1644511149
transform 1 0 51612 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_554
timestamp 1644511149
transform 1 0 52072 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_561
timestamp 1644511149
transform 1 0 52716 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_573
timestamp 1644511149
transform 1 0 53820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_585
timestamp 1644511149
transform 1 0 54924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_599
timestamp 1644511149
transform 1 0 56212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_611
timestamp 1644511149
transform 1 0 57316 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_615
timestamp 1644511149
transform 1 0 57684 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_617
timestamp 1644511149
transform 1 0 57868 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_629
timestamp 1644511149
transform 1 0 58972 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_641
timestamp 1644511149
transform 1 0 60076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_649
timestamp 1644511149
transform 1 0 60812 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_661
timestamp 1644511149
transform 1 0 61916 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_669
timestamp 1644511149
transform 1 0 62652 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_673
timestamp 1644511149
transform 1 0 63020 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_689
timestamp 1644511149
transform 1 0 64492 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 1644511149
transform 1 0 65228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_713
timestamp 1644511149
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_725
timestamp 1644511149
transform 1 0 67804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_729
timestamp 1644511149
transform 1 0 68172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_734
timestamp 1644511149
transform 1 0 68632 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_746
timestamp 1644511149
transform 1 0 69736 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_754
timestamp 1644511149
transform 1 0 70472 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_757
timestamp 1644511149
transform 1 0 70748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_769
timestamp 1644511149
transform 1 0 71852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_781
timestamp 1644511149
transform 1 0 72956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_785
timestamp 1644511149
transform 1 0 73324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_797
timestamp 1644511149
transform 1 0 74428 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_809
timestamp 1644511149
transform 1 0 75532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_813
timestamp 1644511149
transform 1 0 75900 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_819
timestamp 1644511149
transform 1 0 76452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_830
timestamp 1644511149
transform 1 0 77464 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_838
timestamp 1644511149
transform 1 0 78200 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_841
timestamp 1644511149
transform 1 0 78476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_853
timestamp 1644511149
transform 1 0 79580 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_865
timestamp 1644511149
transform 1 0 80684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_869
timestamp 1644511149
transform 1 0 81052 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_881
timestamp 1644511149
transform 1 0 82156 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_893
timestamp 1644511149
transform 1 0 83260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_897
timestamp 1644511149
transform 1 0 83628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_909
timestamp 1644511149
transform 1 0 84732 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_914
timestamp 1644511149
transform 1 0 85192 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_922
timestamp 1644511149
transform 1 0 85928 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_925
timestamp 1644511149
transform 1 0 86204 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_937
timestamp 1644511149
transform 1 0 87308 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_949
timestamp 1644511149
transform 1 0 88412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_953
timestamp 1644511149
transform 1 0 88780 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_965
timestamp 1644511149
transform 1 0 89884 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_977
timestamp 1644511149
transform 1 0 90988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_981
timestamp 1644511149
transform 1 0 91356 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_993
timestamp 1644511149
transform 1 0 92460 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_999
timestamp 1644511149
transform 1 0 93012 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1004
timestamp 1644511149
transform 1 0 93472 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1009
timestamp 1644511149
transform 1 0 93932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1021
timestamp 1644511149
transform 1 0 95036 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1033
timestamp 1644511149
transform 1 0 96140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1037
timestamp 1644511149
transform 1 0 96508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1049
timestamp 1644511149
transform 1 0 97612 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1061
timestamp 1644511149
transform 1 0 98716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1065
timestamp 1644511149
transform 1 0 99084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1077
timestamp 1644511149
transform 1 0 100188 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1089
timestamp 1644511149
transform 1 0 101292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1093
timestamp 1644511149
transform 1 0 101660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1105
timestamp 1644511149
transform 1 0 102764 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1117
timestamp 1644511149
transform 1 0 103868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1121
timestamp 1644511149
transform 1 0 104236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1133
timestamp 1644511149
transform 1 0 105340 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1145
timestamp 1644511149
transform 1 0 106444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1149
timestamp 1644511149
transform 1 0 106812 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1161
timestamp 1644511149
transform 1 0 107916 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1173
timestamp 1644511149
transform 1 0 109020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1177
timestamp 1644511149
transform 1 0 109388 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1184
timestamp 1644511149
transform 1 0 110032 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_1196
timestamp 1644511149
transform 1 0 111136 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1205
timestamp 1644511149
transform 1 0 111964 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1217
timestamp 1644511149
transform 1 0 113068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1229
timestamp 1644511149
transform 1 0 114172 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1233
timestamp 1644511149
transform 1 0 114540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1245
timestamp 1644511149
transform 1 0 115644 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1257
timestamp 1644511149
transform 1 0 116748 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1261
timestamp 1644511149
transform 1 0 117116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1267
timestamp 1644511149
transform 1 0 117668 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1273
timestamp 1644511149
transform 1 0 118220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  Flash_106 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3220 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_107
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_108
timestamp 1644511149
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_109
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_110
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_111
timestamp 1644511149
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_112
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_113
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_114
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_115
timestamp 1644511149
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_116
timestamp 1644511149
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_117
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_118
timestamp 1644511149
transform 1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_119
timestamp 1644511149
transform 1 0 39560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_120
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_121
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_122
timestamp 1644511149
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_123
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_124
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_125
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_126
timestamp 1644511149
transform 1 0 33764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_127
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_128
timestamp 1644511149
transform 1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_129
timestamp 1644511149
transform 1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_130
timestamp 1644511149
transform 1 0 46000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_131
timestamp 1644511149
transform 1 0 48392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_132
timestamp 1644511149
transform 1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_133
timestamp 1644511149
transform 1 0 53544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_134
timestamp 1644511149
transform 1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_135
timestamp 1644511149
transform 1 0 57960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_136
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_137
timestamp 1644511149
transform 1 0 63848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_138
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_139
timestamp 1644511149
transform 1 0 69276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_140
timestamp 1644511149
transform 1 0 70748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_141
timestamp 1644511149
transform 1 0 72404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_142
timestamp 1644511149
transform 1 0 75072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_143
timestamp 1644511149
transform 1 0 77188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_144
timestamp 1644511149
transform 1 0 79856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_145
timestamp 1644511149
transform 1 0 81972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_146
timestamp 1644511149
transform 1 0 84364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_147
timestamp 1644511149
transform 1 0 88780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_148
timestamp 1644511149
transform 1 0 89148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_149
timestamp 1644511149
transform 1 0 93012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_150
timestamp 1644511149
transform 1 0 94576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_151
timestamp 1644511149
transform 1 0 96416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_152
timestamp 1644511149
transform 1 0 35144 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_153
timestamp 1644511149
transform 1 0 10304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_154
timestamp 1644511149
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_155
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_156
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_157
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_158
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Flash_159
timestamp 1644511149
transform 1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 75440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1644511149
transform -1 0 69368 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_2
timestamp 1644511149
transform 1 0 65044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_3
timestamp 1644511149
transform 1 0 86480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_4
timestamp 1644511149
transform 1 0 22816 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_5
timestamp 1644511149
transform -1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_6
timestamp 1644511149
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_7
timestamp 1644511149
transform -1 0 14628 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_8
timestamp 1644511149
transform -1 0 37996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_9
timestamp 1644511149
transform -1 0 40480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_10
timestamp 1644511149
transform 1 0 35880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_11
timestamp 1644511149
transform 1 0 100096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_12
timestamp 1644511149
transform 1 0 117484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_13
timestamp 1644511149
transform 1 0 117484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_14
timestamp 1644511149
transform 1 0 117484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_15
timestamp 1644511149
transform 1 0 112792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_16
timestamp 1644511149
transform 1 0 117484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_17
timestamp 1644511149
transform 1 0 117484 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_18
timestamp 1644511149
transform -1 0 87032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_19
timestamp 1644511149
transform -1 0 86664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_20
timestamp 1644511149
transform -1 0 89148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_21
timestamp 1644511149
transform -1 0 2116 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_22
timestamp 1644511149
transform -1 0 2484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_23
timestamp 1644511149
transform -1 0 2852 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_24
timestamp 1644511149
transform -1 0 3220 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_25
timestamp 1644511149
transform 1 0 117484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_26
timestamp 1644511149
transform -1 0 89608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_27
timestamp 1644511149
transform -1 0 89240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_28
timestamp 1644511149
transform -1 0 91724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_29
timestamp 1644511149
transform -1 0 88872 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_30
timestamp 1644511149
transform -1 0 2116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_31
timestamp 1644511149
transform -1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_32
timestamp 1644511149
transform -1 0 2852 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_33
timestamp 1644511149
transform -1 0 3220 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_34
timestamp 1644511149
transform -1 0 3588 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_35
timestamp 1644511149
transform 1 0 32476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_36
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_37
timestamp 1644511149
transform 1 0 102212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_38
timestamp 1644511149
transform 1 0 101200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_39
timestamp 1644511149
transform 1 0 117484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_40
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_41
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_42
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_43
timestamp 1644511149
transform 1 0 103316 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_44
timestamp 1644511149
transform 1 0 103684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_45
timestamp 1644511149
transform 1 0 104420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_46
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 118864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 118864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 118864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 118864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 118864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 118864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 118864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 118864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 118864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 118864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 118864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 118864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 118864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 118864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 118864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 118864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 118864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 118864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 118864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 118864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 118864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 118864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 118864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 118864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 118864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 118864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 118864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 118864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 118864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 118864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 118864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 118864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 118864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 118864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 118864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 118864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 118864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 118864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 118864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 118864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 118864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 118864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 118864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 118864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 118864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 118864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 118864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 118864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 118864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 118864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 118864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 118864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 118864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 118864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 118864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 118864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 118864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 118864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 118864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 118864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 118864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 118864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 118864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 118864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 118864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 88688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 93840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 98992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 104144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 109296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 114448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 91264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 96416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 101568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 106720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 111872 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 117024 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 88688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 93840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 98992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 104144 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 109296 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 114448 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 91264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 96416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 101568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 106720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 111872 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 117024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 88688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 93840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 98992 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 104144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 109296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 114448 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 91264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 96416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 101568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 106720 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 111872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 117024 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 88688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 93840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 98992 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 104144 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 109296 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 114448 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 80960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 86112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 91264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 96416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 101568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 106720 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 111872 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 117024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 83536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 88688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 93840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 98992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 104144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 109296 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 114448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 80960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 86112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 91264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 96416 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 101568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 106720 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 111872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 117024 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 83536 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 88688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 93840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 98992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 104144 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 109296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 114448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 80960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 86112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 91264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 96416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 101568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 106720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 111872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 117024 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 83536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 88688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 93840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 98992 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 104144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 109296 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 114448 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 80960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 86112 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 91264 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 96416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 101568 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 106720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 111872 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 117024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 83536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 88688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 93840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 98992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 104144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 109296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 114448 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 80960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 86112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 91264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 96416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 101568 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 106720 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 111872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 117024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 83536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 88688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 93840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 98992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 104144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 109296 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 114448 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 80960 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 86112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 91264 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 96416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 101568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 106720 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 111872 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 117024 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 83536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 88688 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 93840 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 98992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 104144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 109296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 114448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 80960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 86112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 91264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 96416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 101568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 106720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 111872 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 117024 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 83536 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 88688 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 93840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 98992 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 104144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 109296 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 114448 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 80960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 86112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 91264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 96416 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 101568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 106720 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 111872 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 117024 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 83536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 88688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 93840 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 98992 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 104144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 109296 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 114448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 80960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 86112 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 91264 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 96416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 101568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 106720 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 111872 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 117024 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 83536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 88688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 93840 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 98992 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 104144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 109296 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 114448 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 80960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 86112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 91264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 96416 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 101568 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 106720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 111872 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 117024 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 83536 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 88688 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 93840 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 98992 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 104144 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 109296 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 114448 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 80960 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 86112 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 91264 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 96416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 101568 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 106720 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 111872 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 117024 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 83536 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 88688 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 93840 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 98992 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 104144 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 109296 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 114448 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 80960 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 86112 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 91264 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 96416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 101568 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 106720 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 111872 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 117024 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 83536 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 88688 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 93840 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 98992 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 104144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 109296 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 114448 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 80960 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 86112 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 91264 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 96416 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 101568 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 106720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 111872 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 117024 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1644511149
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1644511149
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1644511149
transform 1 0 83536 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1644511149
transform 1 0 88688 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1644511149
transform 1 0 93840 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1644511149
transform 1 0 98992 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1644511149
transform 1 0 104144 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1644511149
transform 1 0 109296 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1644511149
transform 1 0 114448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1644511149
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1644511149
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1644511149
transform 1 0 80960 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1644511149
transform 1 0 86112 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1644511149
transform 1 0 91264 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1644511149
transform 1 0 96416 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1644511149
transform 1 0 101568 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1644511149
transform 1 0 106720 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1644511149
transform 1 0 111872 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1644511149
transform 1 0 117024 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1644511149
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1644511149
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1644511149
transform 1 0 83536 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1644511149
transform 1 0 88688 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1644511149
transform 1 0 93840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1644511149
transform 1 0 98992 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1644511149
transform 1 0 104144 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1644511149
transform 1 0 109296 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1644511149
transform 1 0 114448 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1644511149
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1644511149
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1644511149
transform 1 0 80960 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1644511149
transform 1 0 86112 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1644511149
transform 1 0 91264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1644511149
transform 1 0 96416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1644511149
transform 1 0 101568 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1644511149
transform 1 0 106720 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1644511149
transform 1 0 111872 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1644511149
transform 1 0 117024 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1644511149
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1644511149
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1644511149
transform 1 0 83536 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1644511149
transform 1 0 88688 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1644511149
transform 1 0 93840 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1644511149
transform 1 0 98992 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1644511149
transform 1 0 104144 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1644511149
transform 1 0 109296 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1644511149
transform 1 0 114448 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1644511149
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1644511149
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1644511149
transform 1 0 80960 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1644511149
transform 1 0 86112 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1644511149
transform 1 0 91264 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1644511149
transform 1 0 96416 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1644511149
transform 1 0 101568 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1644511149
transform 1 0 106720 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1644511149
transform 1 0 111872 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1644511149
transform 1 0 117024 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1644511149
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1644511149
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1644511149
transform 1 0 83536 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1644511149
transform 1 0 88688 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1644511149
transform 1 0 93840 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1644511149
transform 1 0 98992 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1644511149
transform 1 0 104144 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1644511149
transform 1 0 109296 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1644511149
transform 1 0 114448 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1644511149
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1644511149
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1644511149
transform 1 0 80960 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1644511149
transform 1 0 86112 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1644511149
transform 1 0 91264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1644511149
transform 1 0 96416 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1644511149
transform 1 0 101568 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1644511149
transform 1 0 106720 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1644511149
transform 1 0 111872 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1644511149
transform 1 0 117024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1644511149
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1644511149
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1644511149
transform 1 0 83536 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1644511149
transform 1 0 88688 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1644511149
transform 1 0 93840 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1644511149
transform 1 0 98992 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1644511149
transform 1 0 104144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1644511149
transform 1 0 109296 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1644511149
transform 1 0 114448 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1644511149
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1644511149
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1644511149
transform 1 0 80960 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1644511149
transform 1 0 86112 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1644511149
transform 1 0 91264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1644511149
transform 1 0 96416 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1644511149
transform 1 0 101568 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1644511149
transform 1 0 106720 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1644511149
transform 1 0 111872 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1644511149
transform 1 0 117024 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1644511149
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1644511149
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1644511149
transform 1 0 83536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1644511149
transform 1 0 88688 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1644511149
transform 1 0 93840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1644511149
transform 1 0 98992 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1644511149
transform 1 0 104144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1644511149
transform 1 0 109296 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1644511149
transform 1 0 114448 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1644511149
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1644511149
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1644511149
transform 1 0 62928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1644511149
transform 1 0 68080 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1644511149
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1644511149
transform 1 0 73232 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1644511149
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1644511149
transform 1 0 78384 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1644511149
transform 1 0 80960 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1644511149
transform 1 0 83536 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1644511149
transform 1 0 86112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1644511149
transform 1 0 88688 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1644511149
transform 1 0 91264 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1644511149
transform 1 0 93840 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1644511149
transform 1 0 96416 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1644511149
transform 1 0 98992 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1644511149
transform 1 0 101568 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1644511149
transform 1 0 104144 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1644511149
transform 1 0 106720 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1644511149
transform 1 0 109296 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1644511149
transform 1 0 111872 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1644511149
transform 1 0 114448 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1644511149
transform 1 0 117024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _116_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 93932 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _117_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 93932 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _118_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 73784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _119_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 73600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _120_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 70656 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _121_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 93932 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _122_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 76452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _123_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 91724 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _124_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 111964 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _125_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 83536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _126_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 83628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _127_
timestamp 1644511149
transform 1 0 70564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _128_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _129_
timestamp 1644511149
transform 1 0 34960 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _130_
timestamp 1644511149
transform 1 0 36248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _131_
timestamp 1644511149
transform 1 0 39836 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1644511149
transform 1 0 46276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _133_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _134_
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _136_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _137_
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _138_
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _139_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _140_
timestamp 1644511149
transform 1 0 43148 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _141_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _142_
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _143_
timestamp 1644511149
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _144_
timestamp 1644511149
transform 1 0 47380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _145_
timestamp 1644511149
transform 1 0 59064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _146_
timestamp 1644511149
transform 1 0 43332 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _147_
timestamp 1644511149
transform 1 0 45356 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _148_
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _149_
timestamp 1644511149
transform 1 0 50508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1644511149
transform 1 0 51980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _151_
timestamp 1644511149
transform 1 0 55752 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _152_
timestamp 1644511149
transform 1 0 57224 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _153_
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _154_
timestamp 1644511149
transform 1 0 52440 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _155_
timestamp 1644511149
transform 1 0 52900 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _156_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 53360 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _157_
timestamp 1644511149
transform 1 0 56396 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _158_
timestamp 1644511149
transform 1 0 59432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _159_
timestamp 1644511149
transform 1 0 56580 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _160_
timestamp 1644511149
transform 1 0 55936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _161_
timestamp 1644511149
transform 1 0 69276 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _162_
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _163_
timestamp 1644511149
transform 1 0 64032 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _164_
timestamp 1644511149
transform 1 0 61548 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _165_
timestamp 1644511149
transform 1 0 61088 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _166_
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _167_
timestamp 1644511149
transform 1 0 66148 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _168_
timestamp 1644511149
transform 1 0 66424 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _169_
timestamp 1644511149
transform 1 0 65964 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _170_
timestamp 1644511149
transform 1 0 68448 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _171_
timestamp 1644511149
transform 1 0 67712 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _172_
timestamp 1644511149
transform 1 0 79672 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _173_
timestamp 1644511149
transform 1 0 73324 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _174_
timestamp 1644511149
transform 1 0 74336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _175_
timestamp 1644511149
transform 1 0 74520 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _176_
timestamp 1644511149
transform 1 0 75900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _177_
timestamp 1644511149
transform 1 0 77004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _178_
timestamp 1644511149
transform 1 0 78476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _179_
timestamp 1644511149
transform 1 0 81880 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1644511149
transform 1 0 85192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _181_
timestamp 1644511149
transform 1 0 82708 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1644511149
transform 1 0 86572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1644511149
transform 1 0 90988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _184_
timestamp 1644511149
transform 1 0 91356 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _185_
timestamp 1644511149
transform 1 0 92276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 1644511149
transform 1 0 89148 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _187_
timestamp 1644511149
transform 1 0 90068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1644511149
transform 1 0 87768 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _189_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 87216 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _190_
timestamp 1644511149
transform 1 0 90436 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _191_
timestamp 1644511149
transform 1 0 91908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 1644511149
transform 1 0 92184 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _193_
timestamp 1644511149
transform 1 0 89792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _194_
timestamp 1644511149
transform 1 0 96508 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _195_
timestamp 1644511149
transform 1 0 97060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 1644511149
transform 1 0 97336 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _197_
timestamp 1644511149
transform 1 0 98716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _199_
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _200_
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1644511149
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1644511149
transform 1 0 38364 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _203_
timestamp 1644511149
transform 1 0 37536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _204_
timestamp 1644511149
transform 1 0 72312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 1644511149
transform 1 0 19688 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1644511149
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1644511149
transform 1 0 22724 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _209_
timestamp 1644511149
transform 1 0 28152 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _211_
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _212_
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _213_
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _214_
timestamp 1644511149
transform 1 0 62100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _215_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 100188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _216_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 100004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1644511149
transform 1 0 104880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _218_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 100924 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1644511149
transform 1 0 104236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _220_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 104512 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1644511149
transform 1 0 100096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _222_
timestamp 1644511149
transform 1 0 97152 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _223_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 100280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _224_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 101660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _225_
timestamp 1644511149
transform 1 0 97244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _226_
timestamp 1644511149
transform 1 0 52532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _227_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50416 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1644511149
transform 1 0 49312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1644511149
transform 1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1644511149
transform 1 0 39192 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1644511149
transform 1 0 38548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1644511149
transform 1 0 17112 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1644511149
transform 1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _237_
timestamp 1644511149
transform 1 0 53544 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1644511149
transform 1 0 28244 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1644511149
transform 1 0 70012 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1644511149
transform 1 0 68540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1644511149
transform 1 0 63940 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _244_
timestamp 1644511149
transform 1 0 75808 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1644511149
transform 1 0 73416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _246_
timestamp 1644511149
transform 1 0 76636 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1644511149
transform 1 0 75808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _248_
timestamp 1644511149
transform 1 0 77280 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1644511149
transform 1 0 65596 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1644511149
transform 1 0 66792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1644511149
transform 1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1644511149
transform 1 0 74152 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1644511149
transform 1 0 73508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1644511149
transform 1 0 65412 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1644511149
transform 1 0 64216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1644511149
transform 1 0 107272 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1644511149
transform 1 0 107180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _259_
timestamp 1644511149
transform 1 0 97796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1644511149
transform 1 0 109388 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1644511149
transform 1 0 108284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1644511149
transform 1 0 111964 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1644511149
transform 1 0 111136 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _264_
timestamp 1644511149
transform 1 0 111044 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 1644511149
transform 1 0 113344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1644511149
transform 1 0 100372 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _267_
timestamp 1644511149
transform 1 0 100740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1644511149
transform 1 0 86848 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _269_
timestamp 1644511149
transform 1 0 86020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1644511149
transform 1 0 91540 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1644511149
transform 1 0 90344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1644511149
transform 1 0 96600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _273_
timestamp 1644511149
transform 1 0 94944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _274_ PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 104604 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _275_
timestamp 1644511149
transform 1 0 106444 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _276_
timestamp 1644511149
transform 1 0 96692 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _277_
timestamp 1644511149
transform 1 0 102304 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _278_
timestamp 1644511149
transform 1 0 48576 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _279_
timestamp 1644511149
transform 1 0 9568 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _280_
timestamp 1644511149
transform 1 0 38548 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _281_
timestamp 1644511149
transform 1 0 17020 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _282_
timestamp 1644511149
transform 1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _283_
timestamp 1644511149
transform 1 0 27508 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _284_
timestamp 1644511149
transform 1 0 67804 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _285_
timestamp 1644511149
transform 1 0 61640 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1644511149
transform 1 0 72680 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1644511149
transform 1 0 75900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1644511149
transform 1 0 68356 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp 1644511149
transform 1 0 69368 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _290_
timestamp 1644511149
transform 1 0 73508 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _291_
timestamp 1644511149
transform 1 0 63572 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp 1644511149
transform 1 0 107088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _293_
timestamp 1644511149
transform 1 0 107272 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _294_
timestamp 1644511149
transform 1 0 110676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _295_
timestamp 1644511149
transform 1 0 111504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _296_
timestamp 1644511149
transform 1 0 99084 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _297_
timestamp 1644511149
transform 1 0 86204 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _298_
timestamp 1644511149
transform 1 0 89424 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _299_
timestamp 1644511149
transform 1 0 93932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1644511149
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _355_
timestamp 1644511149
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 46828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 49404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 54556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 59616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 64492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 67252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 69920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 71576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 73968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 76360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 79212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 81236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 83628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 86020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 89424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 90988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 93932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 95588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 98164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 34776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 45172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 117668 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 117668 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1644511149
transform 1 0 76544 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input38
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 108468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 110584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 117852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 111964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 110860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input44
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 93104 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1644511149
transform 1 0 115552 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1644511149
transform 1 0 51704 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input49
timestamp 1644511149
transform 1 0 117208 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1644511149
transform 1 0 117668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 68264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  input55 PDKs/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1644511149
transform 1 0 117852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1644511149
transform 1 0 117852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input58
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 117852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 117852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 99544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 117852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 117852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 117852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 107548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 117852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 84824 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 47564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 113160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 114540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 114816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 117116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 117852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 117852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 117852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 117852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 101660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 109664 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 117852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 102764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 104236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 55844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 64124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 105156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 117852 0 -1 5440
box -38 -48 406 592
<< labels >>
rlabel metal2 s 2042 39200 2098 40000 6 flash_csb
port 0 nsew signal tristate
rlabel metal2 s 6090 39200 6146 40000 6 flash_io0_read
port 1 nsew signal input
rlabel metal2 s 10230 39200 10286 40000 6 flash_io0_we
port 2 nsew signal tristate
rlabel metal2 s 14370 39200 14426 40000 6 flash_io0_write
port 3 nsew signal tristate
rlabel metal2 s 18510 39200 18566 40000 6 flash_io1_read
port 4 nsew signal input
rlabel metal2 s 22650 39200 22706 40000 6 flash_io1_we
port 5 nsew signal tristate
rlabel metal2 s 26790 39200 26846 40000 6 flash_io1_write
port 6 nsew signal tristate
rlabel metal2 s 30930 39200 30986 40000 6 flash_sck
port 7 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 sram_addr0[0]
port 8 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 sram_addr0[1]
port 9 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 sram_addr0[2]
port 10 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 sram_addr0[3]
port 11 nsew signal tristate
rlabel metal2 s 23570 0 23626 800 6 sram_addr0[4]
port 12 nsew signal tristate
rlabel metal2 s 27526 0 27582 800 6 sram_addr0[5]
port 13 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 sram_addr0[6]
port 14 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 sram_addr0[7]
port 15 nsew signal tristate
rlabel metal2 s 39486 0 39542 800 6 sram_addr0[8]
port 16 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 sram_addr1[0]
port 17 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 sram_addr1[1]
port 18 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 sram_addr1[2]
port 19 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 sram_addr1[3]
port 20 nsew signal tristate
rlabel metal2 s 24306 0 24362 800 6 sram_addr1[4]
port 21 nsew signal tristate
rlabel metal2 s 28354 0 28410 800 6 sram_addr1[5]
port 22 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 sram_addr1[6]
port 23 nsew signal tristate
rlabel metal2 s 36358 0 36414 800 6 sram_addr1[7]
port 24 nsew signal tristate
rlabel metal2 s 40314 0 40370 800 6 sram_addr1[8]
port 25 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 sram_clk0
port 26 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 sram_clk1
port 27 nsew signal tristate
rlabel metal2 s 1950 0 2006 800 6 sram_csb0
port 28 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 sram_csb1
port 29 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 sram_din0[0]
port 30 nsew signal tristate
rlabel metal2 s 45926 0 45982 800 6 sram_din0[10]
port 31 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 sram_din0[11]
port 32 nsew signal tristate
rlabel metal2 s 50710 0 50766 800 6 sram_din0[12]
port 33 nsew signal tristate
rlabel metal2 s 53102 0 53158 800 6 sram_din0[13]
port 34 nsew signal tristate
rlabel metal2 s 55494 0 55550 800 6 sram_din0[14]
port 35 nsew signal tristate
rlabel metal2 s 57886 0 57942 800 6 sram_din0[15]
port 36 nsew signal tristate
rlabel metal2 s 60370 0 60426 800 6 sram_din0[16]
port 37 nsew signal tristate
rlabel metal2 s 62762 0 62818 800 6 sram_din0[17]
port 38 nsew signal tristate
rlabel metal2 s 65154 0 65210 800 6 sram_din0[18]
port 39 nsew signal tristate
rlabel metal2 s 67546 0 67602 800 6 sram_din0[19]
port 40 nsew signal tristate
rlabel metal2 s 10782 0 10838 800 6 sram_din0[1]
port 41 nsew signal tristate
rlabel metal2 s 69938 0 69994 800 6 sram_din0[20]
port 42 nsew signal tristate
rlabel metal2 s 72330 0 72386 800 6 sram_din0[21]
port 43 nsew signal tristate
rlabel metal2 s 74722 0 74778 800 6 sram_din0[22]
port 44 nsew signal tristate
rlabel metal2 s 77114 0 77170 800 6 sram_din0[23]
port 45 nsew signal tristate
rlabel metal2 s 79506 0 79562 800 6 sram_din0[24]
port 46 nsew signal tristate
rlabel metal2 s 81898 0 81954 800 6 sram_din0[25]
port 47 nsew signal tristate
rlabel metal2 s 84290 0 84346 800 6 sram_din0[26]
port 48 nsew signal tristate
rlabel metal2 s 86682 0 86738 800 6 sram_din0[27]
port 49 nsew signal tristate
rlabel metal2 s 89074 0 89130 800 6 sram_din0[28]
port 50 nsew signal tristate
rlabel metal2 s 91558 0 91614 800 6 sram_din0[29]
port 51 nsew signal tristate
rlabel metal2 s 15566 0 15622 800 6 sram_din0[2]
port 52 nsew signal tristate
rlabel metal2 s 93950 0 94006 800 6 sram_din0[30]
port 53 nsew signal tristate
rlabel metal2 s 96342 0 96398 800 6 sram_din0[31]
port 54 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 sram_din0[3]
port 55 nsew signal tristate
rlabel metal2 s 25134 0 25190 800 6 sram_din0[4]
port 56 nsew signal tristate
rlabel metal2 s 29090 0 29146 800 6 sram_din0[5]
port 57 nsew signal tristate
rlabel metal2 s 33138 0 33194 800 6 sram_din0[6]
port 58 nsew signal tristate
rlabel metal2 s 37094 0 37150 800 6 sram_din0[7]
port 59 nsew signal tristate
rlabel metal2 s 41142 0 41198 800 6 sram_din0[8]
port 60 nsew signal tristate
rlabel metal2 s 43534 0 43590 800 6 sram_din0[9]
port 61 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 sram_dout0[0]
port 62 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 sram_dout0[10]
port 63 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 sram_dout0[11]
port 64 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 sram_dout0[12]
port 65 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 sram_dout0[13]
port 66 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 sram_dout0[14]
port 67 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 sram_dout0[15]
port 68 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 sram_dout0[16]
port 69 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 sram_dout0[17]
port 70 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 sram_dout0[18]
port 71 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 sram_dout0[19]
port 72 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 sram_dout0[1]
port 73 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 sram_dout0[20]
port 74 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 sram_dout0[21]
port 75 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 sram_dout0[22]
port 76 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 sram_dout0[23]
port 77 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 sram_dout0[24]
port 78 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 sram_dout0[25]
port 79 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 sram_dout0[26]
port 80 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 sram_dout0[27]
port 81 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 sram_dout0[28]
port 82 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 sram_dout0[29]
port 83 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 sram_dout0[2]
port 84 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 sram_dout0[30]
port 85 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 sram_dout0[31]
port 86 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 sram_dout0[3]
port 87 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 sram_dout0[4]
port 88 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 sram_dout0[5]
port 89 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 sram_dout0[6]
port 90 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 sram_dout0[7]
port 91 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 sram_dout0[8]
port 92 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 sram_dout0[9]
port 93 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 sram_dout1[0]
port 94 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 sram_dout1[10]
port 95 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 sram_dout1[11]
port 96 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 sram_dout1[12]
port 97 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 sram_dout1[13]
port 98 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 sram_dout1[14]
port 99 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 sram_dout1[15]
port 100 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 sram_dout1[16]
port 101 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 sram_dout1[17]
port 102 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 sram_dout1[18]
port 103 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 sram_dout1[19]
port 104 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 sram_dout1[1]
port 105 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 sram_dout1[20]
port 106 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 sram_dout1[21]
port 107 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 sram_dout1[22]
port 108 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 sram_dout1[23]
port 109 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 sram_dout1[24]
port 110 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 sram_dout1[25]
port 111 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 sram_dout1[26]
port 112 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 sram_dout1[27]
port 113 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 sram_dout1[28]
port 114 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 sram_dout1[29]
port 115 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 sram_dout1[2]
port 116 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 sram_dout1[30]
port 117 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 sram_dout1[31]
port 118 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 sram_dout1[3]
port 119 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 sram_dout1[4]
port 120 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 sram_dout1[5]
port 121 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 sram_dout1[6]
port 122 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 sram_dout1[7]
port 123 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 sram_dout1[8]
port 124 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 sram_dout1[9]
port 125 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 sram_web0
port 126 nsew signal tristate
rlabel metal2 s 8298 0 8354 800 6 sram_wmask0[0]
port 127 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 sram_wmask0[1]
port 128 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 sram_wmask0[2]
port 129 nsew signal tristate
rlabel metal2 s 22742 0 22798 800 6 sram_wmask0[3]
port 130 nsew signal tristate
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 132 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 132 nsew ground bidirectional
rlabel metal3 s 119200 688 120000 808 6 wb_ack_o
port 133 nsew signal tristate
rlabel metal2 s 98734 0 98790 800 6 wb_adr_i[0]
port 134 nsew signal input
rlabel metal3 s 119200 17824 120000 17944 6 wb_adr_i[10]
port 135 nsew signal input
rlabel metal3 s 119200 20680 120000 20800 6 wb_adr_i[11]
port 136 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[12]
port 137 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wb_adr_i[13]
port 138 nsew signal input
rlabel metal2 s 76470 39200 76526 40000 6 wb_adr_i[14]
port 139 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 wb_adr_i[15]
port 140 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wb_adr_i[16]
port 141 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 wb_adr_i[17]
port 142 nsew signal input
rlabel metal3 s 119200 29248 120000 29368 6 wb_adr_i[18]
port 143 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 wb_adr_i[19]
port 144 nsew signal input
rlabel metal3 s 119200 9256 120000 9376 6 wb_adr_i[1]
port 145 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 wb_adr_i[20]
port 146 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 wb_adr_i[21]
port 147 nsew signal input
rlabel metal2 s 93030 39200 93086 40000 6 wb_adr_i[22]
port 148 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 wb_adr_i[23]
port 149 nsew signal input
rlabel metal2 s 51630 39200 51686 40000 6 wb_adr_i[2]
port 150 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wb_adr_i[3]
port 151 nsew signal input
rlabel metal3 s 119200 12112 120000 12232 6 wb_adr_i[4]
port 152 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 wb_adr_i[5]
port 153 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wb_adr_i[6]
port 154 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wb_adr_i[7]
port 155 nsew signal input
rlabel metal3 s 119200 14968 120000 15088 6 wb_adr_i[8]
port 156 nsew signal input
rlabel metal2 s 68190 39200 68246 40000 6 wb_adr_i[9]
port 157 nsew signal input
rlabel metal3 s 0 824 800 944 6 wb_clk_i
port 158 nsew signal input
rlabel metal3 s 119200 2048 120000 2168 6 wb_cyc_i
port 159 nsew signal input
rlabel metal2 s 43350 39200 43406 40000 6 wb_data_i[0]
port 160 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wb_data_i[10]
port 161 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wb_data_i[11]
port 162 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 wb_data_i[12]
port 163 nsew signal input
rlabel metal3 s 119200 24896 120000 25016 6 wb_data_i[13]
port 164 nsew signal input
rlabel metal2 s 80610 39200 80666 40000 6 wb_data_i[14]
port 165 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wb_data_i[15]
port 166 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 wb_data_i[16]
port 167 nsew signal input
rlabel metal3 s 119200 27752 120000 27872 6 wb_data_i[17]
port 168 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 wb_data_i[18]
port 169 nsew signal input
rlabel metal3 s 119200 30608 120000 30728 6 wb_data_i[19]
port 170 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wb_data_i[1]
port 171 nsew signal input
rlabel metal2 s 88890 39200 88946 40000 6 wb_data_i[20]
port 172 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 wb_data_i[21]
port 173 nsew signal input
rlabel metal2 s 97170 39200 97226 40000 6 wb_data_i[22]
port 174 nsew signal input
rlabel metal3 s 119200 32104 120000 32224 6 wb_data_i[23]
port 175 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 wb_data_i[24]
port 176 nsew signal input
rlabel metal2 s 101310 39200 101366 40000 6 wb_data_i[25]
port 177 nsew signal input
rlabel metal2 s 105450 39200 105506 40000 6 wb_data_i[26]
port 178 nsew signal input
rlabel metal3 s 119200 36320 120000 36440 6 wb_data_i[27]
port 179 nsew signal input
rlabel metal3 s 119200 37816 120000 37936 6 wb_data_i[28]
port 180 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wb_data_i[29]
port 181 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wb_data_i[2]
port 182 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 wb_data_i[30]
port 183 nsew signal input
rlabel metal2 s 113730 39200 113786 40000 6 wb_data_i[31]
port 184 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 wb_data_i[3]
port 185 nsew signal input
rlabel metal3 s 119200 13472 120000 13592 6 wb_data_i[4]
port 186 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 wb_data_i[5]
port 187 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_data_i[6]
port 188 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wb_data_i[7]
port 189 nsew signal input
rlabel metal3 s 119200 16328 120000 16448 6 wb_data_i[8]
port 190 nsew signal input
rlabel metal2 s 72330 39200 72386 40000 6 wb_data_i[9]
port 191 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wb_data_o[0]
port 192 nsew signal tristate
rlabel metal3 s 119200 19184 120000 19304 6 wb_data_o[10]
port 193 nsew signal tristate
rlabel metal3 s 119200 22040 120000 22160 6 wb_data_o[11]
port 194 nsew signal tristate
rlabel metal3 s 119200 23536 120000 23656 6 wb_data_o[12]
port 195 nsew signal tristate
rlabel metal2 s 107474 0 107530 800 6 wb_data_o[13]
port 196 nsew signal tristate
rlabel metal3 s 0 24080 800 24200 6 wb_data_o[14]
port 197 nsew signal tristate
rlabel metal3 s 119200 26392 120000 26512 6 wb_data_o[15]
port 198 nsew signal tristate
rlabel metal3 s 0 29112 800 29232 6 wb_data_o[16]
port 199 nsew signal tristate
rlabel metal2 s 84750 39200 84806 40000 6 wb_data_o[17]
port 200 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wb_data_o[18]
port 201 nsew signal tristate
rlabel metal3 s 0 34144 800 34264 6 wb_data_o[19]
port 202 nsew signal tristate
rlabel metal2 s 47490 39200 47546 40000 6 wb_data_o[1]
port 203 nsew signal tristate
rlabel metal2 s 112350 0 112406 800 6 wb_data_o[20]
port 204 nsew signal tristate
rlabel metal2 s 113914 0 113970 800 6 wb_data_o[21]
port 205 nsew signal tristate
rlabel metal2 s 114742 0 114798 800 6 wb_data_o[22]
port 206 nsew signal tristate
rlabel metal2 s 116306 0 116362 800 6 wb_data_o[23]
port 207 nsew signal tristate
rlabel metal2 s 117870 0 117926 800 6 wb_data_o[24]
port 208 nsew signal tristate
rlabel metal3 s 119200 33464 120000 33584 6 wb_data_o[25]
port 209 nsew signal tristate
rlabel metal3 s 119200 34960 120000 35080 6 wb_data_o[26]
port 210 nsew signal tristate
rlabel metal3 s 0 37408 800 37528 6 wb_data_o[27]
port 211 nsew signal tristate
rlabel metal3 s 119200 39176 120000 39296 6 wb_data_o[28]
port 212 nsew signal tristate
rlabel metal3 s 0 39040 800 39160 6 wb_data_o[29]
port 213 nsew signal tristate
rlabel metal2 s 100298 0 100354 800 6 wb_data_o[2]
port 214 nsew signal tristate
rlabel metal2 s 109590 39200 109646 40000 6 wb_data_o[30]
port 215 nsew signal tristate
rlabel metal2 s 117870 39200 117926 40000 6 wb_data_o[31]
port 216 nsew signal tristate
rlabel metal3 s 0 9120 800 9240 6 wb_data_o[3]
port 217 nsew signal tristate
rlabel metal2 s 102690 0 102746 800 6 wb_data_o[4]
port 218 nsew signal tristate
rlabel metal2 s 103518 0 103574 800 6 wb_data_o[5]
port 219 nsew signal tristate
rlabel metal2 s 55770 39200 55826 40000 6 wb_data_o[6]
port 220 nsew signal tristate
rlabel metal2 s 59910 39200 59966 40000 6 wb_data_o[7]
port 221 nsew signal tristate
rlabel metal2 s 64050 39200 64106 40000 6 wb_data_o[8]
port 222 nsew signal tristate
rlabel metal2 s 105082 0 105138 800 6 wb_data_o[9]
port 223 nsew signal tristate
rlabel metal2 s 35070 39200 35126 40000 6 wb_error_o
port 224 nsew signal tristate
rlabel metal3 s 119200 3544 120000 3664 6 wb_rst_i
port 225 nsew signal input
rlabel metal3 s 119200 7760 120000 7880 6 wb_sel_i[0]
port 226 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_sel_i[1]
port 227 nsew signal input
rlabel metal3 s 119200 10616 120000 10736 6 wb_sel_i[2]
port 228 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 wb_sel_i[3]
port 229 nsew signal input
rlabel metal3 s 119200 4904 120000 5024 6 wb_stall_o
port 230 nsew signal tristate
rlabel metal2 s 39210 39200 39266 40000 6 wb_stb_i
port 231 nsew signal input
rlabel metal3 s 119200 6400 120000 6520 6 wb_we_i
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120000 40000
<< end >>
